PK   �rUB/  �c     cirkitFile.json�\[o۸�+���
x�ȼ�m{���=�>āAIT#ԑ|d�i��_R�/�d��p��P/R�ř��ͅ#�߂Z}��"�j����uQ����^�٣:��f��(M��X��}p��~��+��ê*u�,���L�Jd8d<�C�$�q�)�k%(����=��)�(Km��8�h�áJ�qJ�F��<�3`fS�BG�Lqc�`�1�]��%�P�c ?��h)�O�8�E��)l�,Li�R��8�A<djvbjs�B�Dk�,ա�	5A,��8O�S����@�c	5�u25�j�k�k�k���w�<��*&'%U'�Oo���=w�{����v�耩O9��� ���#BZ��25%���N~y:�9�5 ��2��̧ӱt�l�q��KZ-�x`	~C�k���R�)�J�s��E�EJ�EJ�E��"E�A�'��A/�_L;1	%"�0gy" b� ��0��a܂X*iӢ8��D$��A1������Kb\�~R.�k5�A
�䖮����Z+�_�k�zޙ\����ZQ�_�ka�A�E��֊�l�/�֍j4��+����X���/R�)̋�EJ�EJ�E��"E�A�'��A/�_�����c?�~0����A1�b�)�A1��b�.���8�}p)�Ź�K��/�e\��}q.��R.�s��r�/��+�����-��KpςǢ���j�R�-LUXՙ���[��o��$�f,�j'fv����?e�S��C"�?1�s��g�8l�'�v~:r�T0A����A���g�T�M�[��!���������e�
��d|V����*�CR� 3�?��s�lU ���wƟ����-p$ kx<��0p����eT�m�r׻�}��<�5�7Em�/�}t�v�!�б:S0�:��c � �K(����PPD�	H���;Q��7�A��CQڶ鏶T�ȱ<m�CH�(&P�m���ny¹SQ��~8w�ݜйM���n��ܸws/���w9��O�ҹ��Y��|�:����,؋)2[��k[����}zخ�B���-kA����͟}�HZ���RbKڞ�ڣ��ؒcK�-��r�V�� ���.^4V�0�@h��ew'�4�("2DY��3J�t�T�1�Y��6�q�tB��Ї��$T8��q�2���Z1��tV*uc����G0��H��kq<,�7�L>�����@_��.� Зb`w�!�-:�M�q� }�v:��wco�.U���������+�ncԷCx<D�!2���~���x?�mQ��"��ʒJ���H^-�ź�ۉMhK��!爅,O�P�qe(N�\��"���o��J���-B]˃����Λ6�N�yw���/U�̵o�wu��uS�6�=�J�ffV�n��hVZ��َ΂�j���^��b1�훲0�����������j��fp��źH�zw�����΂�Ƭ�l؃*7�J�M��s*��uy�R��oJ��g9�uѴ?@p]s#!x����ZHƺ���Zu_AFSe��s��Pka̜3
�(�,Mejt3UE�ʴ�q�-fAU�|��,ج̥��ӥ�zbI����n�� x��F���
����1���h�&��;c=��MٍE=��➯�MFc��#�|u|��f9"=EiGNɁ�D�!�Kz�r&�01>�ܘlz}t�{4A7��t��������d&�&Q7�"vb��������y�l������� _��L �7�ۚ�gǵe*�7Es���6�Ǭ�w�3bB�z� 2ÒY�u�E�a�K)�Q���bn�[�u�46��Ei�F(��q�s:�8D�8��:A�\R��u̅]���uqC�Q܂i�J=����s0w�LLx�	�Q���̨���S���#w�T92�e�+lv#nv����b�&9�i�s�K.���l_�ٸg]�����r�#�v�ɑ_~�ݏ��	f�����N�~7��x@����Q���S�*z�����g��X��,�ѷ��n!^IWo�����kU-U]4_��]��rp��Ɩ�g14�h��b�b{xW������-��&Q駏u�)��/��J�9��/���}�_���J�ÕOM���M�Ί���Ӻ�G��`w^�*���_zR�np'�W�2��t�ڋjc����C?�Sotn����M��.�MU��87	�$x�I�qa�r		�2�pb�Z�0¹2�8"(?�	N��1�9����zy��̃����/���?�%�)�"a<G"��qI�wm�4�%�q$9���S��d1кbS�숩���܊o�Q7AH���=YsoWe�a�{���xo)i̮�@̆�/ǜ_��-�����]��]����B?�i�J�-�o��R�<��o�4fs%Tmܬ|��C��η�t�����lE���OՌ�W��[U�	N��oe}���m,���ف�m�]۫7����	a�m��f�[�c���H�6pΑ�}��N 6w��ds�C�6�j6�vO����_�j�h`�!Ѯ��<��	+�dʧ��eS>�L��@�[iʔ��IO���8\��E�[>aA=Fu��oXg������P�'����N��a\w#���d�6�٩�b��g���!�9Mx������jk�#p`:BNT���jdv\�����d�x�M��� ���[�s{��s��Ꞡ�S+U�T�C����c��J��d��U�9�����gl��J<�	C*"��<����D��Zr6��ɦ1����O�Lw�3�<�;�,a���j�`�G�Αl[����u���b�|��Q���\7V��C��ިr���W�����Of��PK   �rU�#��g (t /   images/85cf0215-4010-4105-9e1b-ea712a483bd2.jpg�uT]˲7:���	�N����u�� �-xpww�O��.	���"{�sλ�~߳?�-F�������=�Ǡ�s�� ���� !(  �2ى{��@Z�@   x@A�s��z�6�������-)�P� *�v�6Ƃ�!�G&R
!��/��Ԓ���I٘XY��� =Y���Xx��YIY9�XX! "��o[�	x`�́��?ÿ��4�:ą`��-�{.������rP��%~��7�d�kD�?�������" 
 ���ý@���GDD@B�BEAFF�{���E�OBL�OHHJ�DMJ�@AHH�M������AB�+���������
�������1����a��h((p/@����;zGa`_��# "!CП#��,,����b�xE�*��dO�����@!R�[y�����) 	�5.>�jZ:N.n^>Q1q	I)iU5uM-mS3sK���������Wৠ��а���Ĥ�/)��y��E�%��u��M�-��=�}���LLNM����/���olnm���_\^]���=������4,,,��_P����/�X�^	+�9b���#`����|C�`W>�6vG¡�X�:}v�g����ٿ��_ 
d�`0 !�z��pC�q�+��VŒ�-0�T4�[C{��9�C�N������)G\�-�V����MI��j�pY���y���$���۰����9�)ʕIDE�"c;��]�L�sN�jl)p�Rw��\"3`��`��*�'�h#��o�{��V}%�G)?w��|M�Z�Z�¯_��-p.+���l<�&�-����ih�7�?���{�>`�W��,���ެ��"�0��"t���g6t	����{�m��S�<�o��
7�JGo�r<V��j���c߸�4��t�H�$³�)�kdz���Л��V�g�I�/g�p�tY���t؁j~Ug�Qhi>=�J��ŏ���9���jq��S$WB�$۲�e&`@�v�G�rs�����V���k�����#J���D��.|��� ��+IHp���I�%�*�$og�4�5������DK���Z�~�l�^ކ�z�&.�Si��S�u�2���@�U�����|���L��	��/��B�<��$6��܄x��N����8�!1;��^��K�Wx� :˶���/]&+�,"|l�Cx
f^�2n')ג,����_�p�1�1��m�7���>X@�xr�i=O�_�ό�;0���g%ԸS/}�[�u�r��U�3wgq/1���a�i�2�� �Ӥ�u��t��e��/8I�xf����2D1O� O�;��Uאy���+���9����`����hk��5�?{�#u7�*i$D�ehX�^17����<�~X����?��z�]�yO���Ch�̀v^�{2}�����~��P�t�n6���R��*1�f\Y�]�n��l����p_G�J�m������D�'�yMo��+$N�|�C���~�YG��>DƟQh��2��~��o�Uv��(^�;�NS��Nj}L%H��,�z�@z�^W����;��cFKc��[V����:3���$���~\I��AT�k�0�uz����H9�2j���WNa����K��TVJ�+���_<��$�f[8�q�h�yŧ^���_�Г�q�� ����w�G���w��xe9��-���/S�cyeɄ��%+J皬�JyhP�W%�`�t4(�="VV����ۻ+H���/4��ɇ&�>ۣO��|ϧ����>��CH�`��1ΩQ}�8e�[$,-���Z���rR�`4�^��N��u�+��E������
���/W��eF�X#�n�����4�N
��(S�祮Y����Z�U��-Q)�gf�GV�|Sx	?�����K�hKO�>+r�>P?�)"�*_Y*H[|�>��5
@�x�5Q�d�I/��3r9���e�VC���]+|���V
5�Fʉ���E�?vU��u��e����t�>�f��1U�.�7�S�'�ޫ�/�<���82�#8ܟ��hP	��ո:�����cY���om8务�	;3���]���\M����
T�����-[�CK(?���}k
�O��������N��n�f�r�Ej�u��>0�RX]']Ua���;�~��� ��rRkp��Iͪ7�j1 ��kYX5q7]��(��~Z���f�c�P.M�>f���Ne����ߊM���*[�k��U�i���iI�"�[����=�w�;�a�?Xk��V=���������v�"�J��/`�n�)���u�r�j�dΎ�����Ƣ���s;��ɖ�6g����8���"�W��þ��5���ri���Κq?�X)u����s~{��$��EQtR�;��s���3k�:E�!Lb7�p� �����S�֖�`��֯�z+�B�u����݂6Zs���ܽ�Ĭ��>�}a{`��O�_
1
��N0Cƨ���f�h�������zS����<�8U�A!�J-��S���8����-��L�k�1hڤ0�_�c�@X����`���ro�`&�p����?(��V^~_�I>ʾ(%��(����Ӣ[X}�Z�%>ywF1
��@��F�z8/�j���(ӽ4V��l��K��j�W` �l��$���c��i���)E�{-l����&��prvU1���^w��>�X�>����j�~M�\trA�1�u��X#��^DSQ����.�BS_p/�j|�Q��%m���`][i~��E[E&�񂁘�~�Wt�IW&�`�Ѹ�wc������Ћ}�ㅳ�anaX�W�6˷��$=W׬�(r3��N}�4s�#ga(�!�c,����(��C���_`� ��cmb���u�ק�4 ����.4N&M��0����0{/s?���4���>��N:��;�<�$�	/<���:
WP�ܤѝ�|�cưz͸&��*L��|��Hj��A�>F�T�=���I�U*���k���1�m�"���ȣ���-�z���Y������_�m9���Ĵ�Y߉���:�RKq�.~��RWk�':�(u�z���
d7+)!����;)��Q��s�3qM��m�/{U���X��P��9m��H>A��4����s%�)x�0���7ă6�'\��T���.����|��}��\/�z��� (�ˮ��T�k�g�Ǻ_h���/o��o����{��3�`���RB0��U���$)��V�k1%�N�$�T�x��x����v��ܛ��0W�i����vסw��\�qj"��'�*��*؟���lo����}{����O睑�A�lT-�L��^W�M<�f��)}kIm�JD���k��^Jɾ:���TD0�$3<۴ʻ�RO�p�w?{I��|����l����wS8�_��V2GG�M��	�rS��޸a�m�{�􍙍'�!�*+ΦB���U-H��=�����c��r*����)��+C�x����R2��=1�:�]İr����t�AZ�3y����r7-	Ѣ/S~Fl���s_mAT���}��~X�D�t���z��%��|�����GWҪq��R]j�E���+�C�7)����03%RxD	���2�旅_sL�ח_ت(Gv$F^#�ȓ�h�w#��T$��c��K�派�/����yD����o?�L#?2�Y�}i��~U��$GoV�&|����w{tG�s` UbU���F肫r�9&x��ffV��^�^
���\�{PG,>�ӓ�A�^�4F�o�� ɩ�"ɝ�PJ�?&wĩ�+C���[ɉ�s�s��8�C_#W�3M�h6br84B�*AOg�W�n����A��Cx"	z��-Qnβ���$.+;�%��u\�'��5T��tY��MOm.�'�0�n���]}����2zC�H�Z~ٵ��
ecz�xG��~:����c��7d�3����Sa��v��y
�oB>ñ�ֲ7�M�]\_i�'2_�my���4�Ә��䥃��M��m{��=g���{ޥ�2m;�g���4l��Iʴ�ei^��<����Kmi�*���c*��Wf���E�V����(��G�⏤ȹӅƉwHb��&�2N��y}�3�H��g�g���
���Iӕ�:FD����Ԑ�懛��r�o?qt��v�ks/��6o��홃�ɨ���`.�O�5�Gֽ�)GLZ���s�%�g�k?�gi��@��Λ��[O��؏��[4g�(�:^S�\l�M%_�9��vl�h8Ң(�k&)k[#F���D��[.��v�{�@�ֱ"��^�w�A7�k�w�	3��q�h���T���9��F}˄w�w(����k�l�E�����H��ʌm9��b�g���)[	M�MKK���;���%��ks߾�r~�h�[{�3�������>Z3,m��>�6@J7n�:^��M�_��f��FZ��]}ٔF��o��|ךd��<8�jk��I�~�Z�����wd#@ޕ�	�Z���L>:v�3d��;ȣ7ɏ�B��k������V�-�L]�w���ڕ��s�p�8ij=Ϳ~-u�d�/��=��������3�oLrʣ�(��o��D�⭭OuHg�r�kG�p�-1Xԛ�g覲#���,ʴTjc/Qa��ɐX9Vt$ڬ�~�+E��ZG"s�o��:zP~P�m���Ie���?q��
pa�5��J�M�%�Fj^�-�,�SyU�lrt����J�h��̾�`�|�����b�z�������~����SlD��^�������
@v�c�)�\��ڕ���DS��	r������3@Ix�P�d�5i�.�i��R�̇�B����D�Lbx���q�6@	y�u�xhi}@�����H��vr~ٵa۴���}�t�$@\fG3�yOm�
9�>��x�
���_�S���H-7����8�}+�N�?�{Z2m%/NU��dP��ڻZ��%9y��0�`cב6�u��;�Ba�G`Զ]�����Ӈ)��d*`>"�����|d :E"!�p{,�2�im�Csn�� ��d�o]Pu%u{hv+8?�����d�j-^�c��9,-���N֧(򪤁�[wǨ�Y�r�@����#+�WZ,��Wf��h77��?<*��Sx�E�����vX�v�_&fػ+���ݮ0��_��(�|ݔt'W#��N��I0o�1��?��PC$r��Y3�����:�䢏՘+o��1��w���M��L]$i��g��)B��o�0IJw�	綍����&��x��-����r�1�u~c �z�'b���٬c;-7�ܖ�9�t��Q��M�I��q@���ؑКd��/_����(�ˀ�l��R���L_�
�H;N(yYY�;�pe����M�s4��E��%_p2�A��l�e�7gJ��q�����Fs�(��qײ,��^9JO��(��%V&��E�_	�<��Q��O2T�[�5��������*�L]�[��Q��I������H��V"�p�yE˪[�@2uQA��>^�.�0f���;�4�'��e;~�gT�d{��ͧ:��-����/s�A곻���lℴ#Do�|+�9�Y%�"{'7����9(�'���b%>��G�t����pW���;�k�mղJMsL����ty��дU�.������w�=/��
��<���B�{|F��w!����7��u4;��b���x�^�/�'�Z���pM�^��DW�IT��]�'o^�n�)r�ĭ���yrɊMȏ�{��0�{
�������];����I�T�,�޺�i>gm�Ku�����
���P�҈!o�����5�S�'Jk�R���¢��.ⷫ��R6˗js5��Se��)���"�;$� ��:�F1���Qb_�|u��?U;x�o���V�k�dTT�A��D������(���V�s]D�X9��W�Ĭ���7i
�lf�ǌX$I֯���*���ƋZ2����m�Խ���ڒH O�*S9������c�L-��q_��\X+H]��)kX�/�[�	z��pGMw�si佁u]��;b�LC5��nqi�H~a�c��z��[�����Քocx��ޥ�>�t��k��E�a��k�s�A�z(����˰G(l�p��(�j2}c��-:Zo�l�����O����1��"��V���Q�/����5�kmb���V�x��j�M &\��^�����u[�y˽k%�E&�{6�oC��}'h�*�b�ⲕ�U���` ���zo���_�d�OzN@�컟'�mґ��6*�`���w�̼5F�cF���Y�iacx�ل�Dvu>�K�R��_I!��HSE�"�y�"L��M�_���j��$rLZRT]�E�|����#�w
R�3�ԩ4�dgRg5�nn�������%����>��W��u�ԃ��
f
�%�J�G�۞E�ȁ7�G8��Tf��>λ�-����vu���~^�N��8���a<��	��|g���"�x�ƾ:�=�8E�j5�-F�$|f�V;�djO��]z4}m#�ްp&��TNL�ɚ�G9[�x�V�~�_ئVT@�5������e2c��:�R��D�t�d����A��c��j�f�Sox��K8<9h���`�'b����=��	gs}���3��OI��7I�L�4q�޸5*Z���=�BC��L7=���z3}��ߟp˫#���g�[�fR�o31�Ek)��}���錔iĒ>i��+�K����2lH���$V^�K���Kc�!�a��ͥ%1�E��Q��~<��g �݊��g�K<��=�EQB��Wň�Q�	}�����E��v|?o�4]��;�:`��8��>�m~ˡo10�qє ��R6Nv��){0�wV��'���ڬ�lȝ��#��;��H��t��� K���]�%&2����d��z�o�b�'�P��G������h�
B�.9���O�D^��C����)��_w��G,��<H�p��Ѷ�w�9����#9�,BGy2���r��_حy�k��d�������i�7rz�ä�Ϸ?�RdbWe�Ͱ�v��W�����,�h�w�5���Q�)��1}�ldv�f�UXv��t#4��.B2�D��-�UZ���-gitn��/��a��?�Z��� ?�P*�*[be�:�fCGN@�����p��n��o��Y�� �~B���0�%�7s����N����8�G�[<Q�]?n�M��TR�f���ѳh���%K*&u�։�M����e�F\��f�2�<�H��c�u����A.��/���J��p��R��s�E��YR_+D���.f������CT���/Lx���n}>�m���3����:�/cZobWc	iA��g��~E7+�fҏ_ƠVTdf3U��}#�)�q������r�PM71<ϿH��B1$%�qUN t����Vt���j@����oQ?���guݸGx���3���͘+`` ��(��|�(����[]�P��/��G����{��O�h
V��N�5���_�	�
����I��[��l�F+,�o������E��1�cF��e�<��G���B�;R{�8�u��V(5���sVG4��2b�L�~�b�;>����Lh�-�#9>X�;�����v��P��b�3R�,G��[#����Ey�ʱ�&���:)漺ϊ�v�_�����ٺ�ʭ�J�X]F����	�Mn��}{��A2|9Dyw�{y�Nr3V����1^�.;�U�����b�f����My�ܾ\r���e�m�\Y��.Z~��z@�=�ٝg�����'C~B�(���|7p�����}�G ��c71�hdq���E�0�ot=��~��B!K7v\]K�0&xo7L�K�R�q����!������}j����7v9l㯂�jX�ӵ����M����'|2�f�In}M"�+���s�to���ZQ�"X`��$�F� a=�����	zs�G���A)|vV;��X�U91�Ʋ��b���U.�!wnb'��$��~X��՚�1ڍ�\T�<p�M��/;�ۨ��v����UL�D�0Э%��XӔ�W�V��;?����ܙvWO?f[���׎�=�cgy�����MJTF�j#oݜ?oPL7�~k!EGP��{�f��z�(��
���aou*�.�r\G.豉cw��`9ݼ K�>on�Ʋ"ɱQ7>�⬸���_��L"�6@�\�vZ��J,>�V�0������F:�
kߟ�uy tA�_�0'���&��+����mI���>4�w���T��%nnS	61T��ۤ�2	,���m���J�����do����S�Y�{�@�=�#�TkY�R
$p��mB�-x#g��-�y<��=��#
N�:��?��C�����QOQ�5�:���Kq��S�;eh���R����Q%��k����/?����D�}��g��1Uh������5���� e���i�*~T.������W�K���2�˔�B2�7/�_
W1N�I����r�y:p~2������h��|��oq�7���K�0q�;@-E��s�������Ln��*����;1Qkn��"!�G��R>�_7g�S���.��M�g4�����q���1^��z&�I�Vٛ,G�ՙ�����W��F�[�۩�Pp�$��2{Ou���~#���9B~�� }�|	0^��U����eu�
}la���:�඄"���0Gr�'cz�J��ߓZ&]M����c�oNHB%����S�V�O_Gq���8Zv�o�č>M3BN�]39���$nyO��~` A2Th����Yg!���&�3�=�NR�� 0�T}E6�3_���)� 2D)��Y�*m����ZC}I�<�,�:|ƐxߝT-7l:ʩ�Y��]
��k�*G������Î-Pu�V���wj��x��9	����k�t1�����7�9�,�c$�>�o���#CMt<��}���� �J�wW�֨�'�R��������XR���)�<���8������>t�o�SF���s��S�B'����Qw5jv����>���t~�W�2lRQ�fWj��Z�5_�63;��`s���{�E��l�΁���D��	��+���U��*gK�Mu�v�]�Pw��*O��M��I{xP�4*?����Πdm�
�fxXB��S(6�K����sȗ���+�_��h��Wu:�{ˮr�Yɱ.�Y�`�u$��\�pq��B���=Ne�2g�7���ɬR�v�rE�n�l{U��!�T����~�kTOɀ^�֌�&��5^-CuB�L�V�i
���az�U9[�A����\eT�Ճ�2�DtD=�#�$Kd�B������t������0�V�p��#�����tE��W��	)~�t׸n-t���p5���ލ�`�&N�l>6p_=յ=�h\���j���Rj_�î|�F�/�k�þ_Ϫ�D_T�+O�}w��/T_���2�Ӆn���� ��x�c����]�KhyTE��qp3���Ω��5�M�n��ee�ƽ�	�]��,�+.7</O��ie���wP�e��ҭ�乣�?��D�3M��Ĉ�>���|/�e�U�d�}e.�W����y�wt��f�����-�d8�<�p6܄qF�z���2ԗ�"�{CA�7d�뎉�����+�wm�,^�Aq�S���v���ds<�V�04C��M�"�DS�.�����VZ?@�;����2�zC����1i)��C �0�f��z�8^C���WM�˶o-C�.��-�oԼ:��I%ÐQ����g:&�Q�/ �Ua"u*�D�l���wݞܟ����ĭ;���g����V��g��@��_&�z7o�[��k��o97y��]FN|��8�C��` �=��(?pvh0�)�p�Fy>���~|h��R�mW�M����ӛ�7�(uU���V�k�#�͊G��ܽ��\=i<�	(����-p}�Q����rZz�����;��n^�$�ߺ�Nsn~ޓi!{r��ō���v������G���h���E��d��L�iߡE9�ڈ��v>4�n�͊,K��+;Jj�O|�ۍ[v�F�y��g9����BTL�:���֔z��4���b&��w3�sE�AQ�P�X���s�/G�׹���� 4�ɫ��� k�����%��.ګkj�T�=�U����Sg�|�{4j��#���Tny�F���+���d�޿`��r3!���[��@W�\�܉����X�Y�cX��t���4!�uUо��}H�c�c��T�-�.yk�\Up�a�l�!� Z}�:h�hwϣ�ǉ�]+��M��e�ufB�G�=��i��%NH�(��B?{�e�����)�*TL���H/�
1�j�X6ǐY{�n��)w��h뼴�	:yJ�{Q�῾��e��^�D缤Q��r�݆v�h�gA�0M�v�3n��@��T���v�
�����J����1��Oĵ���������պ`��٦(�կ)�i���3�����+���=8>�I;�R���bk����tl:���0Hq%�n`��O;WX���`���X1a�G��V:����3���B�d�帿���0�"�c�Y�0@���8O�_ٚoy,�x���.�ǋZ+��i���p��l�]�TǣL,bءɑF��Z��l̗I+�G4����E_˅E��ǌ�t�Q�6To}x��=�%4��Y�k<�3���_3l�dC�/_	�(,����k�$�OȀ��U�����B��웲7y�t�z���L��.�?FI�UO$_gR�@���i�$� ���y8�s/�����r��S�,�L�fU�Z�P�\�D��3�ܪ�2�l���}1>��J�I�TߙdoO��Yn�2�c�i���6?F_���1U���O��(�F�!̩�����ՙ��';�G��c_��Vz��?��iƪ"8��#oh�#�4H��:>H�D��OQv��SuIU�g�cJ���%�^��	�}�4e����K{�2�_73uN�ԙʘ�Fѵ������+/|�U����G��	O;�h<`������������b/$�<�Fb��$Z�qR?b�(;oPQ��+D�Ag�_� wN��&D=��8�9�@�f��C���9w:����|3^@��`-s����@J�P�x����\i`�W~ �YV���/1��e���7�d�������5d
��F�ի%D��>}_:��>�L��xYr�S�;�!�����}�揼�(ɵ8f�tj����"x��`�5Έ!�Z�ՍF�_y�՗hV��#�{��E����;���FH���cV�#����k)�]آ?@�J��F��,6�����-�H�Fڟ*�MXd��oI�� xe���Ł���Ι����،��ޖ��ȁ������p02�6s!56� �	��u���L�58�Y�D�,AR^Nf*^
�&^�&���B���|��f.F��6v�|���A�3���􏈋� ���{RQ{'3R&&Fq�9D���9����� O���������d�d�������������`t��s1�`�s��G�������doG��ldl��"@N��a����R����֖�igq7����������������������?ݟ��������3�5��ɿd\�l����0�٘�B�9CFae�����<B<��7q}�.-&@�<*���	Ȕ�/�e����k���n���������m���k���������m��i;g#;�g=���Ą���܄�͔ۘ������Ȕ��ф˜��͜�͘����N �22��O{���B��s���qp1��pp2r��r0�A4��r���s���r��>�O��� 9�ߏ�m�\��l��@v�sUA�f*.F�!b��b��f��e�a�ec��[B����0�U�I{ '55ᓀ(2��2���������|�NfF.�N���6��J���M��M�\�Č\� ���;��O�#'�?��� s��+���OȤ@ΐa=�^�*f�#���gd���	g#73S�&�Fvf����这:#c3#VFsSH�͌Yy��� �h���ml����/����.�FNf��y�D �t�D���O�i��s�4���1F�;���c�����
��������� {���A�����������������ѿ/'fv���;��^���5x��(!-'�';:����� l�\��%EH5��I� �x��L��߿���t5�W6�$㳮���K���� @�B�;'6�`.w�g��� 6S.��u��s�|���3�����|,'UeQ~��%��l������9 �����Z�/l��}������?騐�bf���̇B@��� )`� �p!���(C�E������e�L =� {�0��x���[g����gM(" �b>� �x x������  � _����> x.!����Qf �' h��7�8 �B  w������9��� Ί Ӥ �c ���W��n�f@+� HI�7ݺ���3n�[����'m��#�I[�����@�&������w�21�X8��,��݋�!�#A�	��Jk�� <�?I��0�fW6�W�k!����
�B�:�(]��p������#b@(`h"�~����@
�`�,���@0�����@N7�H�3[�T�kX�=3�a�8�Q6��t��N��X"-��Ц�|���x�\�J��l/�5�%8^�JID,�z�U��9|,6���Pr�'��kC�X{���r�jo+�k�hJ�5?Ck9-$IW;�0�8��5�I�ѥ��O�в��j��wW����-M�+`�=J̯=�୹����K��\��d�wh��1�=�G��K<( ������{�$ۛ���7�m���]�Bfa�j�q��c������M�М����BRӀ`ρ2Gt��_8�����ݳtr�5�x/�^��+hl��gz	��.Q�Qjk�~Ԟ<�B��8���1d?�&ߞ��4g��S�{�i�_U��凲��'�w��c��z��A�\�ؑq�j��#8=ڭ���S��or��@�6[�4Ode�n�oe�t��<�k��"����DO!�5^lbf'���t�%�v����K�d����C����#�+gӝ�~���]�<=������ʭU�#�8
:<}����75�{j�����M�D4�?�3�ӽ�y�wm���-�n���}Ԗnw1F�����#�,"~gf�����b��a�E�9uV,Xq�>�k�1��t\�W�[=�����d�y�� �J��l~��ؕ��P���y�k!��M*ct��7��ԲTc�%A�;���J����Y7��4Z�9�T�'&5�����uFL;�-�_J]#w�'4�~V�6�,�wVvzY�������� '�쌯��&m��e+��y��?��|ѾF̲s�eh��t9V�]���H��.n��U/��f(�|z]�~Doȧ"gJV�Ъ'{.٣��ݯ�&T%�5���W�k�Z9\�P��kmۣ�7$�u�mW�ȡ�e��B����\ٗ܉m���-/�T��퉸S���w1[ZՋ"���Fį^r���T�;u�7�������x*8�d"��dI:nU.Q�u�n�)��Al�F^q�4�K9p�h�5*�i���M���5ÒK���)۞X�f��Rz���ԲF�v̛�������h��!���Ѓ��m���7]Y���5Lz���vN3�Lگj���݊r]8_$����-�������1G^�[��7����2�aw�3��㻤2z7�CxX�7�h�R%C��c��iv�I7��:�G|Vr�:j�C)��dN�<m���9/%E�,�����]�5�:+�/�M�9I��4��]��*�w:g㛛�\�b>�#���Gi;"�mp�ni��*�o��(�mR�J���HY�.$�v���H�W΀F���t'�&W+/�;[���Xi7�)�Ium,�Nt�f[xr�a�Z��t왠N������.wb����b.d��� ��ԙ]��s0��侟 *Rf�Sz~~Ѭ���\l�wG_�Yf/R �]���??)$y�j�� 8e�nZ���'#���˽Ύ�.Ԃ���������UJ������W(O\����Z��Ź#HQ :8cO��s��7+��%�{iS˛i��"�H�M�k����y�بt��J&��*�7�aV�U�I/6��)ڏzhu�oZH@낑71Z�u��iڊ���.��R/�6��e~|�����7N��R��nʊH�X�s&���S?m��57���<�:Ԗ~��y�6gq�����BǍ���w���㌩��{�$�O^how3uf���N˦͛�s�hLk�Z��$����Ɗ˭E�I`&����P�8w�]u�Q�ɬ	�L|�D��界����;N�JU����ׯX)�K��$K$s%��4�0st7l<D�Ò,�k��0�1�t)%.��S�����G�'4�jt��7��i���'|��S[&&�*�~�)/�%�n��a�G`J#�wD�P˓�҆��;�t����U/\�G�:5�;�*Y�-�������e�k�ކ����=1�`W)1�5��
\���,Je�Q�F�%(�D�45l�R
�w((�0u��/]+}@�4�i�i�זx+b�1Z�(�jN�Z�n�)t8bh��aFȦ�"d����1P�uE?�J�|��Tf�-!��au$`1t%�	#�C�B��cCC���p�Id�t�`��H8*d�P��7�s�P�����p<����Æ��\S��e��Xs�-Bv0��Q7�Tu$�M.����u/ �������\��:I*.HE3�i���XV��l��:�� .��
�x�X�z�6���Q�[kGb������5#���ߪB�rW]��^b���}��D�c��AF� �E3�|EN^3>e�Z���V9��e
V,g�O&�A��¢e�2�i�Mo��aU�I�gI�&pѡzg��:�3<o��kc+z$qbmjz��|d�G�h�#�C��+8>�֢����:�`i~�yE������Gii:<��m B~��X��6ӷL��-A���Nl"n�C�z^�>���M�qR�戍'_T]����|�:�t�����$g�A�?��v�%f�˫�-�H�"}%q*�=�X[/y��~q�T�J �c�G�|�,m�9U�4B������.1�s��uf�2�#.G���C5�����Zё��]��j������<�
͊)��ё��&~��s)�41��_����y����b�3�=��>��Ы6��2�4թP���k�y�tsȍt�ƴF�cM��Ő�!���T>H.�y�A�(\g�v�]��Ӈ~3���m,��,$o�� ��ڕg���f��t�M������t��;�;�9��kT}�{n����nWeb�S���p���Mu|[[;����"���������+Eߋt�B^߷q�7p�u�$�S��@�z���������8��c���Z�uޜh�oo^e�2�c5-��ZJ<&�1�eY�^���d�dz�"W����r�/��V���uʡ��3���p\�!��q�Z߭�f�����b�q�Dg�>����<�"��>;���������2�J�C-q?c	q(�.���T�c��<�fͫH�)��9�h0@祭�\�z+Ի�����>
.��[�邵1�{���u�m�T��2��ޱ�/�+{d<z1k90���N�%	K�ɐ+t����±mE��"�"�k�����6�:א	�A:�Ei۟��2��Xj�:��2]{*sSZ���Uq���P�6Y}�-Xe���&F��o�}�X�rH�Q��D��c�M���a$Y#�ԎB�y�
�VLZ�UV����7��#�g5�i�2��8轸H�;�(U)�(�UP�#�T#9석�*_����m�q$y��g����#weȴ�=���+Ly��-�Iq���;}6§d�`��o�4�#R��L���N�A��+� ��k6�p�'(Jt�fJԄ�1��@C�ut����9>,���F� q�����d��4�����g6�� X�m6��_9T���\��;�Vﻝ��D�rL-����Z��o#_�2��4:R:/S�I�X;�N0�ˋ�K�~�Z����1�K�{���P����e���*E%�)�&n���.���ZYE䳠9�3��|~ F3�u��L��ܕ�TH��O�ۙ�����;��mN|�w��+&]�rJ�q+�B�����mb����O_����b_8?�"!}	&u@�C����9����x��o=/�
�$�C�����
d�S��#���X�,��Y�K�9���������+����K��}�-����<+�WZB~d��pw�	�,���l��$S5r��."�OA�*g����S���}�^����v
Y�ʡdw#�
��5߉x3"Q̇�~����y�U$���*�7�YD #F�;��0�� �<�{���*Q��e`ҧv�!]3�Ĩ�"��~��_��	�=�������m�_�)��j^��X\M�|e`9�g���i�U������������ŋ�����;l��ݵ@qw/�����V�7V
���9�"s.�ʜI�$cd��@C1����t��~��$��%:&R&�OMq�?$Tlba���z4[)B���li<�?����-{3�05;ըg�����{"��WN.����ݣ���7`�k�A�wӳ�[���.N��3C�O�M&�%�A�8]����Ϭ�op�����[-���QN>A9��F����R�F�`�A��H��85�fL��8�����$*���r�xz��� �`�@���j������>�M��p�#�M��:jZLTTR��Ppnԋ�w#����y�~�K�,�Q�x��w�t�*}�c�e��^Drӹ����nv��r�^!=��w���Ә�{���'��X(��2�O�+29��K��$�r��������}!X亸��Mm���,-�G���6킝:��+��lE��ÚbQ6C���T*%t%m�`x%�ִڱ(���}�i�p�i���F�j��Y7���[~���z;�uW�(�ȑ@G*�b�}OSUP�C��+���c:��4�G1�0��8���3�R�h����H^.�Q%���ص.Z(��T��_LVB%����6@�-� �ޕ:�<=�ŚK{�?�f¢p�fh���䭡��y+#<��1I�hP�jӅ�v`�vusg�X��.wn����Оp�iy��#�M 
q��k�L HF�ݷ@d���d�<��?dڷ�J2*[6��7��X8��}��g7��������=f	6ˑGyez�ݘJ`J�&a���8�bjyv�0{)��bH��'y�2������̫r��M:�c����{�v�
�r���?���Zu;�x�WnO_���젎^�j`�� P�fd���j�������*�^�s%��Đ�wVJ|����kUe�����;���5r�\������S!�oom�_	��g�>��uNgv�Ԕ��Z2�!)y�p�tO0�l��!!�D*Zz��=�'ϻ��)j��A��*ITҚ��x�A���g�Z�t�J!�]m}U���\��f���g�.���x��寨��K$�C��"���/h�wF:8��Z�Iy�ۡ��-s�(=��.;�tf�/bPGYY�H Q�؈R�!�4�E�])�c�u)��`��Z�
d��
�����M*�T�dx\>ˁ�v{}��N�)�X�Sz!l��u� �.)�a�:܎�V�T��5g��4��Z�~��_EM\&l��{{P��+*4�d�@�9a��[��"���㱹�xB�U�mc�9i�����)��k���d�*�@g��e��R���p�q\�z�VL�M*�b$H!
S/s��0�i�M�RsV%�W���*ɣ͘Y��Z⅛h�) �%��G�A��ɻ�2��q��:O�ꁄ�K �S���<��%[f���Ó����'=�������+��jN�cT���^9�i���V�� �X^�wis�������<-Х=��n�|aO���Hc߰���E1�#cmv����ʌt���W�������Q���JzEJ��0쳙��^�h�ӈ�'����4�u���b�q���y.	>�ri��dU�-֩,�l��}<4e���A""��b����
����_TH���@8���fe h�Z�#�"^X��m�<3��t2�~=��w0F:f|��r��<���;J� �zk@�c�Ts��$`)�~vc�� �s���\�����)j�`Gx���ǩ�b�Y-y�1]�rI�Ṳ��7V6Q�h���bԫ�� �Lf�u��n�
�k����%< 6�A�9�y����k �����~���8vd��o-�w@�~����b��i��?�籯�L��ݪs�x)����� G�Xs�s|�zk^�t��8w��bM,�=19<.n9�\Q!�9�Y,�P����M"�_�g0UM��4�!x��Қ�p&�[q��xf�:��Vx���C��@��	���#���K����z
{g�DN:�&g�7�rYLJ:Q�r�V}˄=�M
����`+j����g�<E!�)�@���B
�8�:H1B��L�	;��(�f�@:<^L_%`*��8�����<����![���C���X�y�7�� GdW�$����"	](ib�=��6�;�h���TT���J����Ņ��Mhe�$& 
 ���m6���F?ДMS��m{�VQXU6F��w��QM���U
��l�$��b>������;����'ZS�������DQ9|�4<����= ��;K�N�0� W���}�>�������±
ƥ��V\6��H�
e�4���f.��/,k45_��<��-��1~rI��5�B�)OE�B��7B8���o���q��jM;��[3�245�X�m���`�3ո�����3������;J\�e�#��慰�\�~"����N���?��L�?�dn��阋U��� ����p?a6ˉ�4H��[��Z���5��a3j�������[�D7L�2à��0wc���5w�h�t�s������>�M��͹�M&�3O�/�7R�:z�E���G�C�o��J)\D�]��V�j��F����8�x�ƋV"�7�L@��ˤ׍��Z�U�w���;\_O��n��l�RF~f�˶`�)�y�qӛ���;�;���z?Q�8�^M�)���6����ܦ���|W㶿z���}E��M�T>B[:E������B_�I���� W�j�7լaC����mH�� �G ��C}f�[�^?�@��a�����M�P�M|�R����C��Χ�+�넛!Qes��lXdp���壏Np�U!c��.��@��MO�99䇼�� ��{	ry���bj�%�Ŝ�)HgL��u�HhV��Wlm�ҏ��������+��.���Ѻ���"�
�pl�
A��� ��w5Ƭ�[s�l�Nۛ�=�V*��K�µA8Տ75���3LO}'7��z�H��R�Ը�dT�L D�����/�YsҚ4��L�Em�H�=�x��k�ߧś.�ϗ����a��B�C��l{=��>P���u>���iR�h1�Y`� qN�r��h��Q�.�e���L �8M׳+E*���2G�3N.�+~��|��N�#�7�Q�x�t�����Aj���D�Ot@��G?�g�鉖}2y�w�M0t1r�P�ׄ����s=��j��)�nW���l��jw��:p���pi�i�d��r�)��ɂv�b����N���k:����C�hf��ำݯ�˂���ދ�Ј�L�o�R�C�cl����q���;�D�ԝ��o��.������� ���2=��J8���Q������B�\Ju͘W2ZD�/k {;T&��1,��Hi^�*�[F���z兛���Z����1����s��Q���h����͝l����k�I��8-� �ZP�r���#e��ע��.g���{	�A0����L~f�>tF�H���� ��֮�04�\=!��{���`��E�^n+I��t�R�5�^�X��_�du
��y��kU��y����HS���,��"@�� ����|�~v#R�=�g�؜����"�~T3=/KK%���ڶ�֗�����'��x쑽��D����Q��-��dd�L7��D�rqH���c�A��2�n�m6y�M��k�-џ݊3�$�(�O����7<ҫ�W���*��U�9�E,.A���A�o��T�K�[�tL'~�qƞ�<���v�s:O,���ġ0��X�[����s�_y+ʮ��4�|����,Ԥ'�����)rS��ە{&�Ǆkct�Hm��r9�&�ɉ2j"���*,c�O��6� b[h�
1[i^�;	�κ��vk}��� �Uu�C¹s��n���-O�|)BU�g)Z0.�JTr;9�ϰҨ�^H���~�����z���Td�w�=53���z�NE��"B���:�x .��_���^O��&u�'
#~ԸR��4FNW)I�t4�Ζ�'�v�CV>dzm-���+�iř2��[���U.����x�
��n�HB`���|q
f|���I� Ť�c�5��ש�G�����a�$��)Z��d�N�廙�I# L�����C��ۈ�h$�
����g	��,����hL�����5]P-�x����<�{��7כ�F�H�5�����K�'ԛ�?_�v�J��^}�ˮ[�W�j3������}P���? �yO�)J�P�䛓�E�HB�)��mAM�V�ڜ�L( b�1\�"����7���W�B����?��Q��ku�q�?pJ܌ӟ�$i�-lm'��G�|T��y���T��i/��l�V�j��6��@�~����Vگ;�$��v����:V���S�T�Z�{����f;����x�{��x�>�����]��i����NB�P��R1�d�U+�+;��`����A�l:�k������_;r�Ngx�i��v��b@>�~��鞍ܳ�h0:Dr?�l	3P�҂��̶��G��|I�;���������A�+��[��.W���GX�3��;`i�s	t}��o��n2�c���F>�[��䷶�i�i�_;ug%�@J4�j��_�i�q��t����K� ���g��wtvQ�)c�,���:���i�}7-�?��jWaUO2�ggZHv��9�+D�
�,�i1�����p����
�����B�3Ϫoq���^yRnuS�m$���>'��(q��Ur8�W
!���j�&�dOA@�B��L &/*�z�F�|�����?��*pJ��9�Z�(�Ml��Ʈ�
=�?���>�Rߞ�E�"��e=���T;����|�εF�S4z�#��:	K,����ov�.X����{��p��=�u��hc��ł}�����W�q�O������Ѷ����b�""5F���|��Z���T
vm�3��w��X���4b����R����O��MZ7�ґ����׊ŗ|ȝ�t�>��z��:����k�O	آ���*��>d��c����9�¢���װ�O�C�)C'�Z�zM0s��A�=�TA�cGkc돜�3gv���S�O�����&��&d�Z��Qx������K�BZ�/�@rcЂjR�T���%���&i���;���"=���	�ߒ�cs����?ݗF�t<��*�凗��a�OA�<�aa6�8�����m_�۞��؋��h�]� ���\�}�s�L��vM�xS�y�CD�Àڌ�b�K\t�y�Ϋ����{5��`y%ِX����. M�<�-�v���d��k24�S�K0MY�2��Y���O$M�oj��i�B��V�5�z_�\Z�7�wE>c������;M>��;)��W�a��.��Q����W�:Ƨ�-�*��s�s۳y�u����d��m}'�奍��. @!!2ė�/� MDXhH@1=ݷ�o.��&&��Vׂ#�*�֖�
�e�[oz}J�K?��&p���a��vv��j���B	�Fq�B���Z�Z	a�U�A�Fu�Q �R��I��C@@#~@�����"��|A��O��ph�T�B	�^�=���'���@���}��&�a`�6��@����M���&�a�_T+� ���B@��p(&`@k��
`� ��ko�F��������3H��/_&�"`H��R��%��=%.�p����%����s�ְO�pa " �PR�o R �7UT� **�����eb_Yhb������EtOu����IEY��a L\i	� ����o&�&�p�������b@���
�y3��(��Sf�/PПO�_��Hh(X4tT2L,l8Rr6NJ\
Vv1.n*j�� �/���A��!>�WlT�oUº�Kl#�xhd	���g'_KGv�ZDv��v�VU|���tVE���t�Fv��v�a��6��q�羅�l��dkg��F�l��
��D�B�.q!/A�#������3�:�D�D�b!;A��cΗ��r�ZU��(�1 �����J%l�L�Qe��^��=�ڪ�����=��<dܗYa�[.��y��k]N��6C�>�����$�����3��!�� �K��Wܐ^�N�	����N&��S�K�m�DϵB�����J���N&_jG��$�K����Q��5�q�Xb�A�.��ܟn����̫���!5'|[�wo�K��9����u�v�г�����I3������m�w��_��]�;��X�������W���=�|#��NiS`!w���wW0�+�����1M����le�!`�����0'�hNh�L���7�.��U��@JD~K>^4���������ШS�U����ы��ç���Gk��ꢖf�䫅ű)7��q~������vq�g��3��VyL��@�_��6Ji���=�4̳�6�n�[���{8���16�tau 2<Y	!,!����R��欹 �)~��pH�5işk�R�;L���%��������)} :;����2�l�95��kw�����FF���Bqu��&[������n{�u
��:ڄ�l*<�:����Z��.?������+^�М�q�܈4��[\e�Bfr�zz�Ո62��������zʿ�8�=)�47<e�=�tJ���>�������SFp���8i���-IL�K���'1D�iޥ} �`x�pA���ʏs�ݸ�)�-Lk��2.��3j�Z�]�d#/mxG�R��)�h�@��Q�)��,��r�y0�@��D��o������z
����_�t��o�پ�a�fW�%5�%״�w���Y�_|��TQ��_�iN�ߧ���*�+o�&�_��خ�i8�xgv���K�������+�������P�ٯ�C��[�fW�U�FwSKx:sO�'c#�K��պF�����jK-��D�S�;�U0f�m�-���I��:=�>${��P.{�K	���D3l�7U�YUGA{R,��5�!�'s�485a�1���i�g�� �ñ�3��ց|6��*SK��4y4���j������ԓL��uw����%�j����p�o?,)k��sI�j
:�?��t���6������^M��!��&���$�E&��O�����:����.tu�ل[����?zPc �IC�mL)fVw��C�e����]<�R��Ķ[#&�3b�r>g�r^2L?� �
_�^�5|���e���!Bvw�#T:6^��pn��`,�!D�ǣEqix�>&��^�1�6��j���B��P<��K[CYHv���L'��+�V:	��V�W�� �'l��T��{�[�o*���g���WqE;ӌa��� �욤�����q���n�a��܆OUA����e����4z�I�/�z�Id�Tx4cT!����p�������M��б�l�ſ�T��z�����ɸGɠ�!Zw��8t�O�X��K�G��M����Dמ������jE�9�ܔ���&����b���������%X�-�ѻ�iձ�� r�J�����js0�&D%���\dىL6���Dn�IXA����p��VuCu�.z�m��~s�E��v��/�trJɑ����~s�~p��̱4�D�?r
<����#/}saɍ�򷴭����;��y�������H��0�KA[t��0��|���[�&��'N�|z��_ �O� ��,e:T�ȝ��K3�0�V�WZ�hn�����W�!��T�""��Wt7m�cm֐V��T����izPU��r!uL݈[NY�f����� |ai�D��z�)s�'����7p�@�!>P�x᭽��0b��l��`4���'K�;����~z���AZ�V��SlYe���$3x�>_�l`E��(����g#�sV��5�\fΨ��'s�]|+�1*���F1:��=�r�0D���&�@,*���C9UhW�0�=�Gd_�[��w_�{�s��Kc��*.��L�z\(1)�$g(���$ؿy���wG�qbq���Wg����RU/Ğ������`vF�kė���Q�h�S���"�_�V�F�܌���W��@�}�U4^U��+�/�u���t�y+�1��8\~�9ė�dכ�"k���<���_{n'ߥ��-�O�m��,�/jH���$|ᛚ�on��<ι�enjr��4�:�t	���\�a����	C�$�,0�xķ�M��yŜ�4�&ķH;ķ\��;$�y���30ˠ$�� ���@���V<ww�Й�xi�r0�_q�˯�o.s���\��C��3��QH?B�1�4B��{�o\�`n��U�{��4Ʊ��Ǳo#IX+�w�=�杠y1�����\�'�f�	?��M"�@n��̝|0c���~rA�v����ߞ%�0���`�a�YmY-
K+iӰ�Q�Y�1�YK+C�Uu���@�!�̄�7��ve�1�12�a�hgE��@6C)��0��BaG����-�Wo�t�@�W�?���l�e����?���.��3.H�0�0�+{dڑ\���ʐnlp��14���e'��p>�a���l8^x�SŗZ&��ڡ,.܍�3�myBP�ۮ�3��7��F χ������1΢����L��R��ch�p�?��^��Ն�͋��F�d��܈�{̝�?0kp]������c�Z��Y����@�#$��-��W=�O�9AS]���]�kw�c"Fb�:�v����y&1h����{�,7�J4��Xj��Fvl�o�)�a����8ŭ9먜�����<oX͚�w�"b*�rS5l�7���xi9UE��䀰�J?�V��d�y�Cw6������۠q��=��!� ?�$2��6q_[��o��g��e,UW���"x�րk
n
3����bTR;8��K����^�Aނǻ���5Z�k��.yZ>��Xޱ7�y�S��>������|)X���B������(ڙ�p+C��n��++�6���&c�t�+Lq��9UEX��Ըi�Q	��0�-�V�͆Cj��5�!�8�ɓ��Zq#���sZ�O����H�s\�]]\���y�c�ycMr���wVRhkF�>���*ү�T��9om���}���"*�o�+��/y��+ȊrO����L�H��6-ݡ��%�����R����Fu�uv���7��!�fH^Fi�#��GU�޳}�QƷ�����m��
It���MI��ᆽXWI�������t��"o.�&��_����o�����1WںW1d�YH����}��|��+~�(�ng���8�*#�6R�"6pgj����M��*�s�諣���v[�>����BjеL���)i�����I�?�|͎���5���-�PX��G:_��~V9�r�}��2��<��%#~�P|�Z|8�p^�4�A���m��}�¨�R�� �.PM�5���v K5���ˋ3j�� u�=� us[���E�p\3��� m�҂=C��R�̬p�'U�doW��-	�t�[�#�y�3�[u��ȼ�N��!
���~0�_jL�U��%�Q�#����f%� �"]�	6���Ր��+C&�7�x�_Ĥ.��H��f�m����eY���g{2���	���9�:	}��m홪����I���i��u��q׹�Y�Ӹ_���`Lf>)<���^����3Q��?���n�� 2���a�v��s]:&�ʬtX/4�$t�s��Y��n�́n�Rtd�%<)vh�@���Z+Z��0�c8I����gwb׏W���7HV+�N�E̾��gb�^�\���F)�a�n�pRx+�͟G#@���c\��~Ɩ� ���Mܫ����c�m���,=���,�pZ\x�\�#���W��0� �~ÿ1���D��'z�	���A�2o���J��.L��дL�м�.�Od�ٙ�ި���"���[����Mk��+1S���8���[t�X8�������FGQԭ�����ǋ?�)a�z:r~5(��΄Tý��}��8�M��̌i�%�r�3u����Þ��v�9�Zf�aG��{t�N�D0[�NoĂ䍨�N&j+h��G�J��\iZ]��mG���ã;�����.CT?���C\��B��X�)�}��q�Ƨ�nKu�s�r����x����b�鍵oA�e�Jx^$�:��$�:��O�U�n��A�Tb��J��l4���c_[�Ir��:��Q�&�t��b�3��"��z��/Q�ØP*�	aґ�������L�l���o,��{�<�7�`-2�_`�?\##�6���=�!�m{�O�����}��>��y�FB"������������s�� &�~2r��HG3ϡ��~����M��v@0�e�me�-���ϖgT�m��m�;&m�g�Z�v�S�q褕<�������[=��H��j�o����{�qE^-�`�w�7�5�'��@�K`7�k�p��3>���P�[c��G�Ⱥ���)�J��Q���2��r7��fw�9��HL���l�&tu��R��٨¦6���6?�&���Z�^.��#�	ͽ�"{�T��J5��e��cz2p������)�4Yq��r�Ϩ������~��s3��k�?��R�+�1ƀ�����K�m�-�q+:�1?5����Y`l��Ҫ뇶��hÁ�vy�C��lR���X���n�7]���y�&�T��Q~����k���3��;Vg_� J9��n���� ��O��������e1e�-$mù��Ί܊��8Km�)�G��!�*���l_*pt��Uww�����S�e�:JsFa�;:[�;��cT􆺛��n��ɴe��umg������dTH ��<f�P�`����S�]�H��\�(�$��V�c�\^JTK%=�x��uSH_��0L��1�Z� ���~�]NGNe���`�o\�LY�.t��Fg�5KW�g��mI��h���8Ñ�ִ������:2=�pW�b���+X-u�;��2Cz_��ls�	��S������{���(���z�a�8�L�m{9
�%Ճ|�O-�X��'s�E���<K�qxc.�>0J���J+��R��S��/W�b�Q�+|����P���:�7����$	�+CZOmt���	,��?��t������S�c��ҮZ�n瘱O�e3X�ܽ|ʋZ.���g����&��G�(c���V�]4���?=�o�$���:�>łJՌ�%pJqu���:�T�'���V����)�gpG�)��8�����o�]$Q1�vٵ:w�}� ��Z=$6���ǍC��SY8��R+�]���~�~�v��<���d`�'�Ƌf٦�ӛ���S�j��-�	Í��.��\��������O�B��M�:��O)ԯ#W����Y�.�ٝ�5�R��jōd�����@θ����XF:;�]���HT��L��������G��8�ݟ��"���y��+��$�5��)�~\կ�S��S�wρ�w{SC[�o=��R���AP;sE�t5�F��M3���IqH��^ֺ��Ǚ����IH<��*s���5o��ъ[��^���>���|8��_@ �k�b�GJ��9�L��/���*p�p�p%a����욢�%��T{�*Jِ����M�3���w��"��۸�bO�oS�9�7���������3�F
r
�0���8�D���/��7�ғ��\4(�䑑7ɢ7����xT�ú:�z*���&����W��_M��~f���Q�=��^�/�v��Յm��u�����/^�N<e-�|��;���D�66$O��9ʌoFi�nXV�Vw����Χ/Z� �C��������uXd�g-�ĺXl�kr���P�.W�O�IM0���|d>�����ְ�e�;�6� �d�z�|�LȢ3΢i�� �95~�3w�{(m�p�H��下�ͅ	>�ޑ�I����a�'��3L�+����8q��&���ٹ��>כnAm�?w�#~.j�K'�����ɝ)̵k����<t�2����jp����	��+�󶲦)v��47Y�C>X�>��SQ�3J�c
�ZXjLdƲ��e�_�55#%H3���ɏq�PG�Ұ��M�ÂoT:Ѕ�d�@KO���@��
���{�����G� G%CՄ��ޫ�V�Wm���c�0Д
Z�0�{�m�fY�h$[����oJ2��%0RM-P&?_��$���v��A�"���]U�s�μ���Y���h���|$����6���@��\t���U����\e3�wя���x/���26l�<+�����͟n�M���w_�KD'6���G�Ow"^�_qv���3@nM[�לb������o���W.t0ϔ�erĺ���w�X��,(�;��+�&��6�+%�IT��͓�+��Z`ʐ�N�f%>���H
	.���i>��H�o�&�c�0/��������7x�3��M�9U�{W%�h)�k��;''�+�E1�!U"��+E�o��G>���#!�&!F�I7W:���$[����4��c��ɯ�ٶ�gw\v�j��y��:7�H������>v�xab�����99?y��,	�C�w��� ����8f��ೢ>���~���T�#�V�ƅ����L������Ȏ��T�X��MET�+ ��v��9�+9w�r��R���'�ä�)��6GZ͇��8Y�e3�J0o�q'�e�7w���B�}Y�� �a��v�x�%BR���8߃b�l\�-< zY���HB���"�ͭ&���	"�k#҂i���<�y�]�Z�neぎ�v���g����'m?I]w���(���/7�θ*#˸,��R$7�p�:߱�(�Ϳzy��*،R�\x�o�|�vy��E�/\����"�+M���(�.xx�y[)c��D5�-5��=)!)&[����lB��O�7����+����F��J"v�\�D9EC�9�����W�/�lj^��gGΖ�=g�|��ު�7�iV}x���T]�9����#��0��vK�_,��;?#�a3��-���܀
tp�w�yz5�k�m��H����G���zc��f�T��ٌ�\�[�9��p��_q�^[+O]�����/<%ik&���q4E��6̩Pgv���;���}��Vg�՟��G�^�N�9y��F_�,,�Ɔ��H��X(�o~6c�Mǁ�1��/�@�ϒ��&��#���OH�ի@Çb;�u;`�M���Q}W�(�{؈���	���M>ǝ3�
�S)@�S\-s��h��A��Q�A�UǔG��2�P��~��$٬���v3�5�O�8lQ?-��.�=8�xag++��U�cp�3�@ŭ���m'Cy��~��ek,��A� H�Gb�d,ٔ=0��Ӧ�Ē�)g���{� z`�_$7xG{{(Sn�o���.z�.�ʽ�	]^�u�\���xb���HK��r�xŚ�ԉau�.*z�G�ʹ�U�aT�-ˡj�3a�������/9K3�� �DBTS8��b"����[�<Rw�;Ql�z��/��]'bu�UU��,�]0�-a���8���}�ˬ^�����j�;$�EF-,�Jl�۸O1+���Q����'��I�����(qX�,�C��wm�n��̍/�QX̗c�$��H�^�3����.�/ԗ-��`�)I%��Cm�!�e����pX�����O�K�h�+�ɬ����lU؆3��6���.ˡ����l����5��:�G��f�B]Je�MN 6��攃dCU+����3K����o�,T��n:mY�������$�ʟ�~u\%�^7T!_����-��֯1�p����t@H�[�����;$�5���a�����$���j2�,����+2�RWӆD.�݌c�^*O����}�e�za��õY��߻'���7Rg�_�S��H�%�� �#�3gĎ
V��F��W�HZ��:Бr�z�t��J"(���2N'���ɚg��aϗ��O��-�1am��HW_#��7-$FV?�4ݠ!tݓ���Z�i>V��w/��r�k_�v�o^.��P�ԅZ��D�6��o��:���f(�������,+��w&ݸ���.��N��PA�"�������eqB��+���	�	}��v�kcL��.C����(��S	p��u}�8^ԿqlW? �Z�J2ѻ��!���G��B�'�6�JzD0�����F=���[}d��:�-�?�AkQP)��u'���*����Ϊ0&��K�F�W�M2o	iC�|�،"c�](2V��_tm�\wN���Xu�ER�j��� ~�2v3�B�)���u3�#1��a�<'Y]�>+A6�S���>?}�L�4e\�^�����Z��&����j���CA��Z��_Ml�Vܣm%�X�f��Yu���Z��6��Gt1͆#����"\��v'E��>����a3�2��b�n��D�Jh�[<���G��h����g� ��*�I&ȕUZ���˭[�6�?�{=�S�;���H��yv�8^��ao�\>/½��*�I��"����\�x���G���Z)�׊���?�a֒��S��W{�pi�#��+���`S'N�R C�J�4i��ׯb���eeLY���L��6�F%����]I���|�:9�$jI�s��bx|�Dy�EyD��^���+�UMټ�����C��"����-
0o�3I�JsֲK�¢�-/�?əҘ^�kɛjJ����-� ����3e}JAXj�?@;�F1�-�
����S���̐�W���j��,���P5x�t�\q�T0ۻ���m:�2�E��JP��d����"� ��q̴(҈\EWNd(�>dH�̻����'u?��˺j��� �%r���5�}��)ک# ��ǄNp7�>�q���r�9��c+=+1��2QC��Y�{��B�U���$˥�Jv*�BI$�����yO|Ì�4������6)3ķ�]J�����������m�K�ޡ�]��PI���[uB	�����"�U�M��+�L��X��+�Ɋ^@��df��g0���⑕-na�Y�f�r��h��Q7CU�v,�A�o8i�\5źd��Y�]}�d1�L�y����_��q/CK�"m���TY&�ȶ�J,��x�q�n#�)\�T�Y�sٽb�����D�a<.�l5�&���'n`5~pq|*U�+?=�e��A��H\�H��"Ѯ�с0���Qu���ye ���ӯ+�ð*�jG��,,=<�2y�;�G�_��|��D�
Ή��) 0g���)�6�T���T��
�e/*T�Q!��*��q�P[�d����.(d�=d8��6�M�����=K}�H7�,e�(�r�c�;)�RF)��O�G.\�W�;����vO�L'�n�AH�Ws=�x�_�-i��g���to�.i��(1S�)(k ���u+�H��|�>�������)!_ub�]]��B�;��x��#�c�}�����D���P��Co*���ƧڈcR�s�Ȉ1���K��)8�9XH1�]c��R(�B&�/�a��aE��)"+j�5�K��@s��|zN|�Y���K%�s�LCRKqa�Ʈ��ި�t(a�~������mi�t!K$�O����iH��z��h�\��}$~�Q�óu��R_��iF�v����RA��g#�q�ժ�=��.c�M�q�D���t��G5ou�2���B�nc��5��SyA�P���r�$e^�8Ͳ�*�e���x�w�d�wޚ�ۀH�C:N|�1ASr�w�t�w�$ul��yN�^�lX�3�ޟ�G���`{]N�������?���iK�JҍU�Fj�@>�S�k�,��;<fx�2u���S�����$,���@T���1�����N�o�jhU��|9�*Z�?UT�%��8���:��ͭ>���n7��#nn�4>�ρ�<��0�T���Ha뤳
��Ȱv���H�G��#P� �yd~W�C{�ͪZN��!�?��G�������Z�y<P�q0\�v�Pd0�-�����l>��*��Vz�&��H�ύ�Me���	�w����0�.���R��Y���*Q����}���S��R(�E�؂��:w5�@�iZ_O�F�sbC��JxbC�,�=��	|d��� 4
�GZ+&�Ȯ�&͍��D�e��u��I�IY�[ �,����n���`iggGP&��-.���"��X�
�(���N�P�n�����C�Q��;�;�H�;�8@B���h��)!��{�?;���~fwfgw?����Y[NI��\�8܂!.�O�m֋����ěcȀ�?`�k�gqؕ�̘z����&�P`�z����R�t���/�+�K�K����G�AE��W)��T)
:g��Hi����3E�h�IZi*��G���N8bl��]��.�����W<�ri���^J�1ʜe]�k1��N_�`���*ˣZ��J4wMX��?]S���?]� ��OH�%w6;P..-I05!-F0��?F�?F)-D0��?��I--�1E�8EM�O��������������́K��R��՘�iێ������ bg \^��bxB��������DJ4�a�e�zIFFF91I��8�D�^$Q��H�$��Q���Ǒ�H�|�~��Cͨ�������H��O����K1�� �_ţ2q������ M* >!!1���DD��xK $�fz �K�n�NI�*�VL�P�m��C�z$buL�)�����W�K��-f������%�ÓŻ{�D 3���R�SC-C�m����	O)fە��E@N���^��j�"��ӚI��M�e�Ԏ��w��I� e��: ��K�����d,;��XD����ka%�YR�d�o>,Iti%,���3�A���^nKB�}����B���ph��\���cQ�"|���0�1,-��ձd��%��b�j{I���9Kڠ��W�g�IW��Q7N�b $�9;)�Yĵ�OG�y̩�4��b^?ŵ�X�e�������7�\:�y��:)�z^����Z�#S�z����U	Ґ3_�������G�sDu���ZK�2��J����"�Ŭ����-�^{�{HRx���c�NHkb�{G�ٓ�@h��ZL7U�
�j{4��`ꓫ�PF��B�W��tgz{c��= �'N��$jR�U����|�Ӆw9wKxF�d�6AƝ,���#����T�������;d�'���j�����mI_X��,�]!.�ר�{?���ю�%+ƶ�����/�|[���C����=y�� ���l\)�+d{��\���_���gY�OX2�k8{��_��Ĳ`Ē����"����̝�x2�t��Qϟ�.	[$�Q���*�(�~ʹ���>��ybG����]�@I�>I�v(I����9�h��FV�Q��p�>g�=W_����~9�#��"ջ	w�g(�,�כjw� �}���lq��ښD�7���r��'�m�8��*��S�
�7��K��Aq8���7�8�f� �g+	�X�U[װ�g��T鬛�yz���.W�M�ς�NXv�����xy�J��j�R։J�h���P)�8�= ��PZ��1�=>�#"�v��͓tl�#� �xC��*u;<��a���P����$��twf"/ú�=Y� ��k��Y�[�����3�^��yx>p�I����ӥ�Xa�3�0Z���r5�M��H�y�=�8Y6�!�w�������D���Wx�܈��1:yʜ�#�/tz���sA-�{ ��tU�����i-r<9?����I\��x��ʳ�#�YS)z'i�rn�L?��8^ۘEÀ�*%v�	�.9�z?te	:@��0[[��m����C�l�pX7g*����Z4����_��}�>=���!"c5jR����W�_DT<�l��z�"�sh>�I�̤nzȳM��_,5�S����c��77۳��r���l�%"n��v���O�����-��~־�`�r�L�zo�=����yo���i%#�@Z����Zu����L�	�r��5�+�5V=z��;}dq. M%��sU���.�ߌ���&�"S崊�z��v�}��VR�o�([�Fݳ伩����>��2�*o?+��d8)��Vì�:�a�A��|sK���U��F�L/YX賓\���%*��I��t&\m��t�vȍt����p:�k�8dS.��7]V��
cV�ޏ��#�!Tf�]a\���"�&��������˘��G���b%N����J�h�mq�e���ra+�0B�����u�V3`<O>�q���o禢�ܑ���v6�a�/��=�l�$IV��	�bY� g��=��KE�����>2�(�њ�~�M	�꺘�u��|;%��[���O[_V9�m0�Ÿ�y4��:�#A����r�)��r~��0ޠ�-���@wM�	�
I���s&<U
S���5Xr�Ϯ|iu�`�#�w�g��Xe��Y��Ҕ�b�I��r�N�˚��Q�9�m���,�ۢ�n	ܥ�	�O��2�����-�u<e��q�[�B��3C��8���Ņ��T|�򖄨-:?np�~L-ۃ��B��(�<ٛĹ�Y�@2�#<��#�09Q�F�A05x>/�o5}��(��upE
r�r��a����tBq��>��=�	{���V�����t�NS�-�}W�-�y��>��ָu-�+��5%���/0�\�y5�h��$-BRh�ˌ��ao&[F� 8��C�N���X \�ǋM �O�z�w?�����NM](Cnuh�}D{v&"�;�|�I���"��Dc����T'`������mU�R�^��t6�J�^ϑ�DҐ���3�)ey�
��#xԹ��)D,C��\0���F�8��Ve�;�������-d�,�N�[%:K�1r��S�yz��Yr����.f��ޯ�N%���cr����`{�ɿ9�������s8ܕ�ً�Q�L�dD��������
5}��S눷��S�C�)�+����q���]�Zc�ܺ��)sOdxٿ�A�s�DC|�2(�DpsZw
瘤K����w�r`�����T����Kǩ
Y���:������E��l-Hk�.�FED��]�X��T5�IZ�.��w�2�4�U�v�ˤ@�pB��)�C#kXl����Z���	B��I2�����A��3{ýW�x*��L�O��b���f�Q�ܵ����ʲ㿤Ϲ�kt�U>��|����<�|��t�5f�?�d��z�Kp}J�uCj�L�m3�?��hU{kZN�t�ц��-�Ȫ�����@U[��U�W��+=uA�z����"��J���_�닍2�:���L��!�3`�A�!��B���Ԋѓr�!c�%|Γm��O� �����w��Ϸ���5&��q��������q�":�w��yAT�L�=�4��0�x����`E��]=+�ns��Hiի'={0!���O��Q{�aFv�X4eS�(��n/��mmw�!������9����nk/
|����]�y:6�8�5�מ�F�馀c�c��ϲ �'|2�3l��fE>��8�P����	�/��(e�u n��f)%��t�X-��+���Y7
[6i8P�b��*���[{��Ɩ�w]�'�瑥QZ�/�:������!�xs��vPCFy]E.�����b�����~e1Kқ�M��N��7�~��
�u����ƕ��V���Iթ?Eb<8:3���o�^��� ��'5��`�����a��A_������"D����\j��!��RW97���r��������-P@�(ʂ��PΛ�b�w�����z�?<�]W�M�W�A� �'N�-$eSWc�k���9����Tٗ���3I�?x �J�}7�V[B���*��@u���\��;kK�8w�5-�]��#�����S��3{��EM��O��N@�w|/+c���rB7h�q՗
�+6�P��$zAw��Ɩ~�O�Jd��#�k��H�"ӑt9���m���n�jV򉏛��tO��B��L<h{��v'��rԑ�${s��h-�Tj�P��]�a�`IK`�cs�k~�Y�h�x��{�Q�ט !PC��B4|�)���o����n�T�]���3�EG?��{@�Fsi�	]_����x����"�b�~$�Z����t���xP��y�����Y�z|G/�2-��V�_5?ī����:G��ԧCh�Dܙ? E�o�!
@�H.�� V��ޥbxfD��T�>��x!:���/�ej�^��G����#�|$_=�N����Ȝ�%�E�����*�����*zMɨ�:I�� >*�Y�9'��w�:[��'����!�t;���)��;�sC�J�_�v�=�vH&z)����L0崬��  ��D�[}�z=+gv8�3Sw����U���,QLȸve�^�xv�P�
S���&g��s�� ��j�hAd�/P���'m#��N�x�ܽF!Bۇc���	er�i���7�6�"Y���(�ĳ�d������Ç�f�,���gǅCd��Ȫ�*��Y��'�{@�IS�wt����]^hs������j���T���e�y��I=#÷�y��|����Ob�9"��g��3RϬ��J�`�3����N_��S����.N�~�N�?ˡ��Gi�{4�Pbҫf��]�*�u�Ro�_�v҈E������y"�w��r:�)��C��'�����7�5Ya:Ws��.��e�[I֜��V��f�Eޭ������[[C~�Fljqd���?V�
�YU綵 $rF���Q�V� r�������������[�B|��.��Ar�	M񇌚�ۄ�P�8�T |��@�����kl��Â�= �8�,��ƭy[���ny�JK�Ǖg�F�d�o��ju�B#+~\ho[��־��M�U6#^��nA��"	c1�li�IT���4�mpNe�d�]2�0n�^ �i��oo�1Ld�(�px��*�+P�/�����Ҟ�,��u(T�rD>�w��3e��3͗ad��-g!�\��ږ�~\�}���G�Wه��N�-���}���ޟ��4��vZ�ۘ�9P�M�k�a�Y��("|B�o�@S��0��,�FQF?Q��#��g,�NG���j̊�F���x@�,w��R7�H�<��Y�(R�6B��&�T�
3�6,(�=* �ӲU�F� ^���v�^�10��%�,K~6<|
�'��(�*��v]?�YW�>|
/wT�	�]?W�b���e�R���P[�a��=嚪�G'��G}4��qp��)�
�N���_V&y�©n�������MB�.f��&Z��*e��B��y��D=dp�H=�n�t/Hϧ�*-���D5���ˈ��BX���.�i�>�0�-����+ܞ�I������Y�J�|�c;�F8�ʢj�*U���-�KA����N��xv��<�ԮǪ���*l#z��R8\��tTYnHGq�W���	��_5:��T�9��[�S����wY�
�"�CK����j��jqۊ��x�_7V��]�-�zſ�nk�[��*ϝA���=�7w�YтU9*f�W�g9���c�BC����
������Ũ���m��6�A�SF��OC9�xN�GxW��/��VF}X"͵�|��-�%��t�7�d�U�6V�v�~v�س%�.
8C�]�uj�8�e�/�4�[�������-S?��W�m�0���Oa��.��;?Q�@|^�J��l��?���a�!���!�9�&�;��c��K�/p�w@�(���~~?�L�d�(*~�s��2�g�UP��|zJ"--�'JÎ|�+.����jW�,����-��T�{�k	f�{���F��`Ur��qn�d�IHU8��R�o��qѺ�}��Y��܂lt�'�fTA5I[��!�'��ՎRp`�%`��Ւ�)I���>�5�o���?g�Al�N	岮�9�Q ���y3����c�A��jt�:e0���F� B�Y^�"9�EQG:��U.N�H�R�{����c��g§:���Ӑ���:pØ��o��Ct���NI\MځM�N����U�eم�;˘����b�Y�.��D?�Ĉ��Z��8��8��*�K��˰bt��p�(n�>�<�G1�k\�W��:^�PJ�m��>B�_���A/���O��)\�9g��J�%�{}�B0��I0�D�!t�D�Z�i�~"��l88�|��7h#[��f�����r��xY}���m�#��������)u^�q�^V�w5�:|c;^�8� ^h���;� ��q<��֦�J3�.�^m�[�r�����Q����{ͳ��h=5� s\��'>�3��������g�J���j<��U��ȧ�9�qus�&�w����}�z��d�F��K=�F�J�lӾǯ�Uf�c2~R�����|�N]IZ�5�1r��h��j��x���� �Ut�hU��r����W�������4&�Z#�~B U�	�rݷ̽K��K���c<���C���=�@=�6�4b�d�S|w�,V��ף���
��$">�H5�J�3_6*���c�>ڝ�6�k�Dd㤰�
��������s}�v;H?j	}�ii@Z�&�T��`���ǥ�s��`��-E�Z�=����J�����].���մ��[�.���Cj��~0
��"%�^�ɘ����9���T&��Ood;+a�[a��\k<��p�n߬�[��mhd�R���j�Ց*��F(�¡:ď�B�"5D�;�q�eR��ʌ�By�4�b(��9&�}�ATC�jQ�u-��!b��/��-�H.�PPw���/k�{�B"��C�����V���{\��SI�X���v���$5���k�j�M�ϛ��prI`���s��_S��g��ݘ��)|�Y��:d�e�>��s�\/�u5��롔$����lPo���L�>�t)�虠��>r7LsG�Vu��\�ue)��H�EO֗i�������7�8I��9��L��Ǆ|�:�W+~GTXX�L�d%|1���i�2*�7;�� @~����#/�_"X�-�HGb���H�<��m��.sɜ�ʩf������hv���ͼ���vzpP��J4���V�y5�pC���]�R#���P^g��[�$q�p�qE�m��HF��o���GBڶL]bڲ�7T��S�i=;��s��2�{�C0Pk}�����R���X�B*����7^L����e�d� �h�_�@��b�|��K�W�`��ʫ��/��4�>�a����|i�9<����?��L?����dU�Ml�b��Ћ�h@���.�u9D�����ʝG)]^: �_�.uǷ;�C�%|=&�4���� �K��<�����N+O�ǡ��iyMv"�|��t.h�go�������� 	���{7�6
�K��eO�	��@���$�;M��G��6Ԙ_��঑E��� ���CC��ȟ��-��xx��HW�Mzb��տ��H�9nD��#=*�i��OE�J�z/X������m��O^U��Ǜ��L��\��7I}�&$C�xE��5�04��Ļ+�����Ld���M����D˼��yz�ןw-�0҉�+l�amf�M)G_w�"Y�Ɯ�tu���-^E���� ��,��b$@	����$Z?<��#a���hL�p�K9�FѱX2~�9?c�PA3�II��fVw;�iT)�L�{�q*v��� ��0�U؏L�����$�d�p��n]���8�0v}�8GY�,�<����a�+%V��&q�P�b��X�]eO��WzL�6s{x�m���d�`����t����C�1�w�bE�g[�E(^�f�r��lk� mk�ŧ���r�,�xu���zr����5Fx7����௉��v���>R�&�خ���)��"�n����Pi� 9%V�f.B��t>�_�lk�6����R��O�rT�R+TԴ;P.W��9�,Z9A�g�������@u��9���aq׃ICr蒲� `���~���e��pP�V�Ԑ�.�K��Ͷv�okm�nV�a�^��z���<?�3��ص�������9W�=@o�o[���ܢ��{��l����d��j@�����&��_N���z�,��P�����^d��,�[�Z�R[H�:��fNpGZ�\(ԁC@�j(��q��[��M0����4U�n�=��{Cb#]�)��VK����M��+�(��Z���]J��� lp�������әc݌�=�qj嗅�T]��I�×�Y��\-|����7���K��fp��#�U.0?rF4&���S�sU�ۭ���yv9�����w9�Yc� �Ė�?F#ǥ�Z3nK��i.K��<h���W����aým1�`eB/�ɐ����q"<E������t��+��$��9��F�)��	���BmH��/My�rXS�p��-m1]�JԖ�*�=`�:5�<;�Q:+�Ѯg
2̾��vU�r�5��:�l�y1oS�[6i��>|�8�,W�[&K��xT!66{
���1����o�Ɵ���OQ��[�>ǯ�4���k���A�Wf.h�ˍ\>�L@%RO|a"a��3����BY|��B����F~��r�q��3�1�=�r6��c7�W�?SX�v�������9z�J�����Y+��cN��5*�[-�*�쯋��>vܜ��3��n�&c���'Oԁ����y֨���I_��}��$j�]'��o}j���l���l���~����L�+e2�`T� M�+]-����DVj�4X�ey9��F�N���X+6#w?�d5�{3c��?aD��`�����8�����]�����L��n�x�c�S��*��^N8B܄�ӃHʁ�r�yUEM���ګ���^l�%�uEY��!��j�C��Ͷ"�������aHX��X��c#|�G͞�.�Px,�L��;��"2�4��B)߰jߐhv�Pі�l���ɋy��!�����?�a2�u]z�o�m&��x�U�K�?���mʡ%�淖�(�W�zF��o����!�w(w����M�ޤ����kO�\�77H^�>���P�������];�)�ݩң����v�.P���+��-��.xE�=�k�g�d8\��lH��$�r��Ty��R���!�rT"4��|�u�����?��oG�1�^��恴�d��5LA��3���v����HEc���z��b2��V�д�������_}uV���f� �GV�+<�v��O
�0�|)�z�����Q2�	���D@H��*E�5�>3͵�f��b�r[��]<�ʨY{f�}jn��m#w!Ck��:̷#Q��P,!T�f�	��k9��j�h~nQl�%ߤ܍��Ȃ�>"����hd>�T����|C�[�DOƠ籡˛Ê��]�t��%��X�;t�L:�K.m<�'B��A��5F���er��K�-HV6Y�r�~q�"�.O���#��0ߌ��ȁLSVj��t1]�2�W�@����"M��Q�z�<�q8��b6,�_dsu�6䕣ʻ�	BPRw�ò#��c�jV��0�y#;���av�z�])�z�\��*��G���ʪf�y�a�r�?��N+��������/1����VǮ'�0�!Qó�/��� ��u7��/���/MR���ج�'�Iڻ߹�����O��wPO��ɻ�e}j,;<	F�R ������+Ğ�ً��m�A�_U�[��-��V����a��c�^&�A�����=s�%]R|�k�b�_j}#�MlT��Sq}Xެ65����abu��%�_���,ܾ���̥�T�ylX{4������%�Vp��q���d�;��>�@Y^?�\�lu`�h��7~w\���pú�Yy��gw/���1�����
��;�Q�
.����]����3����c{��:���723N�n���<��e���f:?5�j��[�C6mj���b>뺜[��<�ƮCz&vr���l�9if\�������l�Iա�����
=bH�kT��-XO��X�'�0nX^��-/�MQ�j�0]�O+���o�1��6��ݤ�^�1]�͉68�?���F����&������zBp�j����Kvo�tg@��F�{��%�l�Z���t����x��O+w�@��ä&�60#B��왕�����~O�ѷ�^� �'Q�\���Ř�l�}R#���5����V]�><<#z����.�	��"7G	�jx:?��7�����x�3�[S:e}��i�I L�h_���������D5bUQjQ����Z7Zz���g�Mv�\�V��v���"�����l�dQ,(�N�D�+��[��`ȱ�L��.�ԩN�Tt�J���{\����i:�m�	~��Qq�*97c3a�ZN��Þů�����W&8������jU�a��/~o.���_ԛ��9�F�^����k0oE�ݦ��vPV=���̐������E4K76�8��,�\�	�
u�~��´C`�Y9�'U|�ʚ&�Q̖�5o����:��!�|45��K��zЛ��[��4,OfRL�e�OQ�:�9iwVN������_E���u�YC�	��Ò>{AO�uD�r��II\�`�z5�a��D��j���� ��R]��6��]�ihc��ǐ��\EIY�Bs�>�5�eY��_mG���� �^7>c���Dȃ���g/ xK>?��(R>Z0D�tO���"����u�L�Ŧ�ܣ�k*�@����k��ij`�-՟p%�+}"��i�΁.�K���Ҟ6C�ŇϜ�M(�ˎ�ҕ�$���lb��C�9��\�����*Lo��-:�uث���G���p=o�jMw�OT7���V)�l�4MM�uA��S�L�M�)1��eu�"�T�����r���d<��p����B͑�@@��S��c�:,�r���h�<�Z�ps]�\��g��b	��o��J�Zʳ�̯W䩛�{W³%��x����N~>N�M�p� �n��ƭc'��|��"zx����"!	�wSH��t���-ʜ����}�z*d�ߚ����8y�>R[����)��"Y-C�/.�R��b����i:'�Me�ᨺ-w��J��P��bh���r�t�E�m�e��� ��ٽB���t8:ҏ"P���S�@��kC[�R��GWҖ��T�E��ݢ:�rK������|5Kļ��مe�V�]��a����l����0�k��Ӵ�˙���W}����ӭ�4�R^54�]�ڿ6�:{��r6W#lhjǪ.qS�k���-�����m��a�� P�ɣ ��a����|�Gdx����|x�#4�m捞nԤ�w� �U�dw�h�X�/��C��z���f9���!���p��0w��k0��g-}R�ư	9���P+jߢ<���3c��!�S���},�|�e�B�j
zF}>A{��{Ԥ���-�u*��=�M����D���j�=���f��a�%D�(��=�O�+&������}�g	��nU���ɭb�ο�m(����Y0�p�y\Ki�"ZI�v�Tho��H�R��Z������U�x�ɺ�sl(C�_���-l��M[~��6���N�;���Y�92J�f[����'�?y��W̎���>�mzƽE�B�����~�I�~��M55�P�`�0_��~�@^��L�� ��e	ՏTl0�ef�G;��-=��lVzʖ�J���P��(�/��{�T�[:�Xw�gZ[��I�HK�qK�5_M���ў��׬��Ϟ�b��u0_���kb�9�Y  ������fP08g��ʿ����r+r�����}5��̱�6���طOP�����&0�Dݯ��|���/S���
�#����D�-b�v�i,�����m��W�k��
�P�1{�6�}�b娀;:��������ᵤ�����+�[LT�V=��6��ɔ6��EO��2���6	&�e����Ӏ9ǚG��*}j�|.�C�٣"O���j^xF�16��f���r�'$�dǐ��${/���{�a��.a&tMY�~��A��^�*#1Q}�K#���^l/U�T�׹��Шz��������P��t7��I�!���rENz�؛[\�Z�K<voý�GD�.���::�������H���֍�͌�o�]`֍l
�2�g�� {6V�T�-�sHa�/��(ya���b�u�T�t��uLp���#�_�I���Q������1\J7<�i�kf,}��.�&�*ޡ��G;ƺ%˾ڵ�\��7-w�y��*�8��8�۾<�����Uc�	YI6�e���A��z��(gN��Grӡ�������|���q��E���@Փ�����ErIRG��r�
e���s��r�(:	SGF���9�O,i�	0�ᱽ>��9F��r����G����@�D�u	"�Z��G1��'�2(oKېH�_��x>�C��b\ջD28*f����mI5���O��x��rB*C�9���35 �MW� NE��O-����a��O��ͭ��NJ��н7vU�A�o���M�4vPx��;�]0���?�c�
78�[L�����M�+Gp���a�34gK�JL��4�ƍw���)7�@�i�v��V����4B��o��z�:[�"��6���S��!�Y)i�C"�X��ɉ< Fg��iT*i���������HE�Q��C�j4��[ۣ�9�J��:*:�|���%VR|C���~Z��87�~2���\�N�IP�wv����MPmg��w�cr�%t�hA���7�x��U�&l�y�M�t#40���f�Y#=������FӢyWټ��AO���2�7	�H��EL*:��Cwn�"�8�çQt��W�7��LQp���6��H����;=�yÁ�6W� �8����p�XqJ�[O��Wy��CH{��2��è�n�E��ZoT������m�LbX�X-�� �
��:2J�1E�e�����j׏���q��+x��j梉͹�'$�w�s�?�.ᶦ1:5}�ƺ�^{�?���2�����}������w�֚�= ���yV�d���J������C���E�[Z;X�P����OOI�e�oFU�I��P�E��y+��d�'\Ơ��;4�B8)a�*�!�L/�)���h��˻�9�zr�D�
5CӦ�ѓ:E6p߸�E���=#�f�.�Gm(�ۭ�$r����X=`��tA�yFˌ��$U:a�H��/�|����C1y�b~i}ZV��g4d}�*;,cv��Y�t��Q��!�QԾ�%V���-I�\5����E���XY��/^��p؜�Q-�U�76	�S64�y	Åx�TD�o��f˷�7�c#��ˠ�_��͔J�����}*z��g�;�'�;8ժ��\fB]�:���10`��!�Q�Ș��a[l��*x����'8����l���o-�ĪI&��.�i����H�+�}c�+e��g㯙�*��O艢,%ć���|ɢ�@,LkRЙ�wޮ�dd������Qg��V��u�sђ��\z�ꐂ"w�
�:|���,�$�$����쫏)SIc�J�U4�M=����{���b��r�_M.P��Ƣj�̶�����sN)k�x�e�tȨ���k+@���	�|/~�ZB�U�� 6�x���¶�{H�ݚ���7S����s��B��@�84�*�]q׼����{0�u��O>��l���mÕ.X�Y�
n�9`��9D'O�Ȗ��j�x�$d���,�e���]Z�����>W�W�%��&,��W�ؾ'��)�8����_��F�F�mSm��ٜ3E���.�����`\.�~Q�������eX���t$OI�ԤC#���!t癑�4�l�1Z�;/ǯ�
���[����Κ����8��n�J���2P
�����U<t*b6�>���0Tt$m�!���P}�����]�$�A��Nr`� �>Fp��M��C��qd9���Swi�H,��ʚ�I��hI��k�܀�n�޻<ӗ���!Q�Ŷ�<Y"b��BI�x���=Ϳ�ޡ^���f'#?��*s�ƞ�\D���*�������K�庩ҤU�J���4���W<}3��64�*��P����Qel�Ok��u�#Ɂ���5Q���Jk��QI�[���j����%�e�/i��Dw����۷�FwO��E�r����G5,��{Lǽ�YjD$�<�"�h���<D�wA��xt�j�7Z�R���k�
�>!
��P߸9��e�Kq��퇚5k��t�Bhϋ�����Ɉ\��V�r���o/Z)��y�{@{^$]贽�I6�T�Xx��%+χ+�r����xf�ET��rh����ʨOu�o-C��1�_�p��d�3Ɖ�W�һᆱ�OߎP���������d�?��E$N����B`�����xT*㉇=Q힅���j[�_ƞ	=�ϸ~|��Zw�)�wM��b��~��5���(ڊ��P���5��Oi*|�ب�������܄�l/�azc��qղ����Rn���e�Y��U<-��3�ә\����``ܦSZ��I�!�����a
�(	�Q���Z��Ϧ{������2��'�x���ٞ�ک��~��N�Oe)@~y�E���`R25x�E�����QO/���J�b��Y��T��qe�Oo�yMͿeqhb�0�E:�[I���\A�����6�+=�PD䁺s*�p5w��緣=�K|�q��3)��R@��GV�:�,X�g�c"�����0���h"E˻�vD���Oi�j?�]�淆3�h~���'.̤r�0&�(�3�#li�O˪��GyMS�X#B���>�F��O���zC�u.G:���r揂�t�ũo9�����W'�(�4�.�:�`h����ף��va����+����E��z���h���6�q����G:��l��YRt��Z�t��!�Fn�χf��7Ҕ��r�����w����P5H[���=����Q��}�:oN�Zr��>"�!���d<1��{�R5�=�W��.�g2�&���T�݉��㙗]>�A��G@p�OAwi��qZ�%L�C��$O>L�k���T���C|y�/���l�&J� ��  ً���#w-Bu��O���CsVT�TA��R⬧�x+&=��F�sG����ſ���e���{Q�5]mU�T�
�#���w��*��)��8���S>�fO���(�̌�"�ȯUg^�����o~�93&<Jm]c�pRk�M6�\��?�@�	~>��L`w�o���G�j���(P+��24�RK9��؟��SM_ΫH�*W�G��:<+�51�jH�ѽ�U��sy���Ms3�_}��"��7˞e<8>�E��W��p/A�B�K@����v,�uE�#��r�ٯ�f���Rk�}�>2�
�~�ݽ���#j��:h��{��R���(���><-7=��d�:����}��������u��&�F/o
��e�&a���<r,I"=��Ȏj�xF���-՘�u������E�'tu3��Wp�g3��kS�q��IE�\��Oe���P���E�%W�wBӒ�]��¿{����nߟ�$M2R~�4����+!-�4�}T�y��#y�዆6Gr�y�+��D��?)�5���%�s�]|s�xG{���~�x\��4�n#;���qVF�1�Ʃ�nÂ�<���n�q���;��tMfU�iS��~���:��)d��&{��yyr�j�1B[�7��^���&U������x�A$l�z�q��A�BM�>3�y�k넥`S�t���R�v�]F� �VB$� Sb�d�1�}��S�$��Q��qѱs�\V�l�qل�y�o�ߙZ�H�'%��TN�᪲���T��Ŭ�Iy}��$���+Do�����'�/��st�Ne~�F����Sr^�>����wB+��V~=̺�1/�|;W���}p&0ɘ��F��.nr2�E?I�@N��d���
�@=��E�++���[���"y\=5崅��)�eޘ(Ǭj����.��b�E�|���&����2��O)c��\ƱG�|Ұ
�.]p��c�n6J��w����H�0�񖲁��i��z�&�Ǽ	S���mH騨P[QJ�p"�8��׀gH�Դ�2�)h�!�3�>J�e��w���Y��s�m���T�ǿ�%�����Z��Rm?x�6�˽�NS�S�   T�Ċ����l��j!�e��̩���k��J�=���h�i��y��.��=�����@*�jٕ�9�����-9���t��"0I}��J	�^R�a�|߯�B&�?'9�iw�d�\4�@q�ȸ��Ԡ�� ��Uػ�CN�x�45�$\KYU5^��	�n�<�"֜��� b@��3�V�;���0�Oά�{$"9jE=�������?��G�	�u��Δ�HrcI֒���Ze��Զ@ Dւi�(A>�����&y�S�L�)(#*��f���b�TR�艠*h�43@��)3ʂ沅'_�8��=̿�h�i �ZJ�O��:oA9<�.(�D�Uf1z�	�|�i���I�@�ր���X^��#ƭ�Ov'H�@��qJ�^j뼉Q����V~���<��V����kj�t���.k��<�,A��5��)��!z 6� T��{�G1X��>kDM-9D�� ���EH�sR� F�5�"�����$�'����X 
#��"B��jdW�����@�Lz���e�KJ��H$���"��3Z�P��}i[���k�5y)�Y��S;{J]���$���'�A���Y��Эrժ��?�'�H)�N���Z^ޘ�+�<!�$'�6�4�P�9��
�B���c0�S*�J|��%4	o�r^�:I��J�V�i*'zNTD+є��A0��Y�F�4�"O�z��)9���.�����F��޷H�)+�1E��֟Z����{�t4ܞ~ш֒�Rb��4���c5���0h��v�M�A�l��4���Q]���b���.B�c�ݺ�g�I�.܏��k4�����:S�V����	�	�ѷ�#.�E�D�,G���)�P	ץ%])H�K��Ε�B(_���#Шާ���$�k4�M(skV���$%'�'x�3�IǢRc��ƔB� ��\%G��m���jw�g3���L'ʛ����?t��U��5�JI15m�gQHINZn�DiHw����t]�X5�*d���T�^�����%�:� JK�=$M o�4�E,R�mJ�+1#zV�4٩iI
�h�%�$x�h��(f�IT��>��E6�V*]�)���Z$tV��zC����CZ�IRG:.RNa4T���}��&�Z���!�zR ����b��؀#\�Oʮ/𵶔/.b5����@��M�Mr�֏��B�~t
�~{R�l��=)w6C��iҿhZxE�^J1J��0T���{b6��}d��@I�z��HX;��Q������Y��eҘ�u���C�I��:������J�O�����a��@z t�$Ed��:G�F�G��2��k^�� 
��hQ�ֻfN��7m�b��N`R�H��V��q�ڶ���Q��V����5�)`{�	�T��Iʿ�(����
Wh�pju���}�.����i�u!d�U�M2�oSGS�◝kZYY���V�h�
ueK����ɈHR���kk��Ck��1�R��•� A_֊.[PJ��u�<��,�k4���<M^�%��A��U�M�� �6�G���/�!՝?�ұ+��ey����� 1�k��~���j��:��5�>��]p�dL՝�q�N�i�T������@9ޘԁW���6���xZm�(=��2'�=-6�k��v̠ ��Oȏ�n�R^����xQ�;����~b�5zL��N���˧�E�r懯���x�2n� ���q&&�	����1��8�XW����� k�17��R�8	�*��y	��H#Uh'�E2�� :g���K��ʕ$4��t��%
�?�ȫ�cm��够�C� m+�1�V
_. k
Jc���q��:�w �v�	��y�~���z�R��<+��ӎ�}�ly*ְ�%�dm�R��V	��[4��B�5�
K,'�@�O*P̒ yW�2�S�5��\j{H?����l�S�j5�N�v'0�ҍg�;WinzWk>�­� V�ev3�Ma�wng0�(��l~�l�A}��}ڸhe�yW�s�������|�aY�	��T��&��.��%M�_j,��-�1yR����;
9GƽaT&���ɎT;�C-J��7��a�)�s�$F���o���!%(6�p�&;�z�o��+
i[���~���N�]�f�X�qb�RJRk��6�'C��r�zH���Q�*ʡ�+��]�1؀s- i��y����Ap~��$��9'��~\��gm)	�֎Aη��KH#Z���jޙw�~�<�Û��{0��)�Kn)���$QpWhh�IRҩ�;���a0k���1j�u���')��|;6����U͒|k��ɂ7�����QYk-@���ՃY��i�f�¾�X� ��Ir�v�ٍ&O��s�Ԓ<@���U�*�+7.��e�wF�<�s��f.�;�|��V��a e�mAԁ��co��Kq�O�mI)qJ�$m��?���Y�@�)9U��ư�G,��[ʩK���� Zh�M6H���n~�ꔐw���B��A'�	��ڐ�i(�
E-z��hFƊ�i�� �:Rď:}����QX�%�T�̔��\Bȷ�NA� 5D�1E�V6��9���ֆ��G:�,R�T��;yՋ!��s��p��
�s��A.�Y�_h�:��҆�3�X����U�`v�R
cMb��h�@��_k��Ѧۃ
|(p�:�(
ܝ��Rs���1���e��
�H?1֒��>��Zu�&�(f#��u���dh3�t
�XKM5V���ΜP�Eu��R�s��ZR�N�ֲ~�(�w�oɍ[]�����#��=���zt�U���1{�N�'$��w�R�$ӣ��&��53�H��|6�vč��\P�=�ֽ�)z��R{�ꨬ)���*�N�V�v�a(ְ.E��m�{R@ x��?����J�J���k��=U�m�# �!)QH9�(��p\ĜN�DJ+�[�y�_B�Vo�D�{���:�����n����#N�VXsjyA' $��:M�&㾬`%jڮ���^S�'z--	�㨮*�M��V��]�B�GZq��)U�3����ՙi�Czw��%=�'HBGҮ;�P2}(�E$�')�e��[��� �cC�V�( �_I�XJ��iS!)P�9��~�p��Y &�	��q®�_/�q;��;��Wi�E��/!\��g�p�t$y�aMt])JR�B�y u�X;���-�n C����9M�Y[�gImm$���4��QW���Z�	RP�k��}�>��:�Md멨�HJ����GݓY�Ƨ6�����:R�#H�⇼5��|����$e��Fo
��U��6�AN�ʏ�E�im�� :s�j��@��wJg�D')�'O�-juJ�O�u<��B�6���t���պ��$�ݥ� .]|�+�JNnuo�[��Oά�7l��;��5y���?
t���>�D�4��Ŝ)�7�S�Ɔ�L�(��|L���;5��I����{��2H�ӂ���6��3�&�_y@R[��Wov ��ұk��î'�'�X��~�yO=|�*IJsF��#ƒ�P�V���J�F��R>i.%�D�W��a�s}a`�R��̝�����u	+�U����%�����֞��./��rjz��t�sI(i.�E8�+Ʋ�Z�+�6Υ����"��4 қAˮ�
=��߭wL��*��5f����8��C�W�+
İ�5ԸBU�ɝi��["�m ��`}�*�^/��,]�ie��>qΧ��uZu��>F�D����dW:�YO�@Ry�(���(�@�_ʠM`���&���<�D�S��Rڨ�+*�B�G|ǗJR�:��Mc7�8����g4� � |�l=2>�����k�؂:�:�^(o�f��e���uZG� �sִ"DQ�fEz�c�D����IYk���;��ml�@��Eb8��n⑪�>t�qՕ�A'�E��T�6��U�4��CJ=u�t��2T4Z���V������*Jȁ�I&h�t��<�	����Gm7��g�U@�deH�&)kD��4��m*b��;҇ҝY쫉-;3Z�]g	S0<����i�uڊ�:F��L��h����|QV�-J�Pu�� ֭�}�-@��T�:�fӰ��2�����,��BB:�S���Kl�/2��� ߕ5��Fm�A�hw۝�RR!)�|k��8�,Y8�+F�	$nzM`�ư�C�[\�d�k�#I���c&%kp���d��>T��xfN\��z*�����c�o�5kkr��vjȑ��� z���K�
�kp�u���Ν���O�\	�Al�g�ޕ�߸t�]$����Ӝ=��i��-�	?]����c� ��LkNp�,�����cQG�x�[�ܹ��z��Z�lէ[��	HP�!#�s� �2�.|b��W^���� H�r���(�)5�!Bs��� I�a���|5�b���<��Ɇ�	�v�E�J@R����Sj��t�\��U�&��]�a<�N��ə$Αp�U�:śj���� q�-�g�^S6����	�<�u�W�������4�HCh��R=:�3��J��yaN��9�k�l��-�^�l���> VT�)#��P���Z��;�'�+�k�m���t��A�&b5� R�(� �VT�ҝ?�?J�ѾD��@
��=R?Jq=������:O3���.��ˌ�S��gÙ2�tO����U��S�D�Ҝ�\%�FD�wF�����HM#���k�$�8?�Si�
G�#�e��z��-�3IߗJ-6����;�O�]`v�r��C�ޏ`�s;���[p6az��BJ��ʎC���HO����φ�}�������T�cƣ�HRu5�s�UȞ�S�s�� ��� I   !1AQ"aq�2�� #B����R��03br$@CS�4��PT`c��� ?�!�v��FG�#�va���L	Y� ���r�t�#�-� �Pi3΍�]�M�ׁ�҅�W�xg�J4�� ��I��;�c��F�P$�w���C]3�i�O٩<�J��� ��� �Ss�B�\u?���]�Ytt�(=�^��z4��:l#U�U����e9D�B�wޑ�P��N�s�Ak���N� ;�!
G�ɬ�Y#u�\|an:���<ФF�O����Gr�4i�"ӛ.���#]g���4I9!����r�ٻ��,���F�����7p�8.�������%�� r�M�I>��<��@��s摴񅐴�O���Yr��]uA��8�6�WgR`A�J���<�M�Qi#}���}�Jxq������������av��������c��0�p�<���_	�ȳ�q��?!�*���{�}��Ѯ� ��� ��'0��v����p�ueҌ:���aT�� K`�� ow�XuN�c���U�Ο:5�0wl鸻R�O濆pW���2ff]�������	�G�3ħ�G:R�k��4:-�7޶����Wv��#���� 4�`�іm��_¸C�&Ճ�Y���1���L�t�~i���d�g>n����!�J^���`�`hp�ot�d�8>�75�xj|S�v�����W=§(�L�'�O���}�|%ߟ�8�b{ �xI1�T�,-�!�3��5�`�u9�.ͼ��a��E�AB�$���U�;�ӆ�p�	O�,G� ����&�kO�G0��rϛ��*�Gp�?��d�tw-ϒ|?���a�L6$q%V���n=쓮Ry�]�M&����Ys��Tz;њ��oQ�vh?ZI��;��C�Jmw7�P�f"i:7����_�Ti����Ќ"L���T΄�}C��;��Bm�pI������ �j ����a����h�:��yR[�u���&�V�7��.Ƒs?=���Hii��T�GG����?�V�gG��]sTҦ�`�*��s�ZT�[����a.?圼��՝�Q�ujoc4�>
���+ٶ�Û.�#T�������A](�f�a���fi�0���Xnb%~�-rY�Vo��v]4�E;&�փ�j[����������Z����?p�����8j�NbvV��,�ۊNppv�WD�X��-�r�*�=G�����ll��i�����i��]"P��^kل@�"�7H᢯d�sk����f�r��J��i��+�=��>�А�J��>
ˤ��A.<ILƨ����B����4�j� ���b�g��1���u6���ax�p����RFi:n����TX*@ӑ���M�O?4��iͰX�7��!�Ϥ�[T�s�n���]׬܎�M�g����.2���2��{�T��� �0���W1{KF]Ɗ��gpk1���5<�F�AK��U�������v��lI^���j!vCa��p}��B���4-ٲu
�ᦩ�������X���I�*8R��$����l�n	nb�܏�=�ӏ�u�4h֒y�J�[�z4ն%uk��I�Tm��Uо���%��� ����p>���	��:��PPmǯ�����N�=��F�z�ov!�W��-/!���8�̢��A��BȝH�0�oksE�tep��9z�.󷵡VfCL��U�(4x���;�Ml�b�hY��N�F��\5+�Y��ԕ�+b-]N6�}ߊ��׽�6
��HK	�B�yuN�!��mV��eJt��2@w�J,uZM��o��A���a�i�]��{Jy����k��W�c_��-pkҤC�.����ZM�hʠA�dqX��Ш���t�x']{[̸�UaزF���Չ�r��]Dj2���H9��ec8�o��tƊ���d�~+��+���Oo��GTh���}*N�XM�E��^�aID������h>��8�K˗Q��fw��� b� �IۈT�o�����:�%iU����C������L~�+ќ�����鯪�<8�2��z'�Ӥ�s�[�	��(�p�c0�?ԃ~���Cw%���h�m"u���k���wg���Y�J{3V0(fʺS��9+�}*�<d�Uh��]�'[�F���z���[Ҍ;m���c6Y�:��v���V�o�O+5��W�|����+��vK�޶W0�mǇ��������F��Qs(�1���Q���&�̫X
q$��t[
x5{�?���HeO�4�Z�6#R�7�G�k(7���!x̎�=�z��E���<d���g�9(;���St�u�"T���6�{1����;
7%��k������3��d���A��}d"I�aͺ�,|�{��j�4�Sx����U�'��]Ul��Y$p׊l{�~���~R�24��q��,4�F��h�*9�hY���	�r
�H�R�u�&�I�p ��';WJ��r��`T�2֍QO��'�����Ti�OU�\"�
䀹�I#�++�ր�#MV(���>��\9��X_T������Q ���
���m&��XݭZ��R �������l�gxi�k궦R�nx+ �}{㓘 j�I׵E�����pO�a$�ǰڢ��H�p��f� -�9��ז�U��4��!��X=�����	� af�!\���.��=�ƦCL|�aټL�^�Цb|gf;B�fkJ�wDs�BZ}�X8�2"`/z+�[�w��д� 3s� ��^���S;�hܼ����C;~+�֮�kN�w��]Vb�~�5��� �Rq��X�?i�)��_�������
�kS3_��o��N��-�YR�<�k
�a���k�Q��	�����K��@DǀV4Kmã+"uW��.Z[p�.#H%��T�5�U��RnC�Dމa�~hL�%oK�-cM�:jZ��%�����`u�-�'E����Ry�O�
~��5�}�Z���d�f�6�����8�]��"��8��Wt��^��ԣP�Gܬp�-�~~�f㢼��B啩�2a�[[��kYQe
M'�� H� qY��*#��:��p+���z|�X���kܨ�<��U
���-�� ��Ǫ{I�j|7V����s�ߏ�D�O�.��m���wQ�p�A������xk�.^���/3c?qT��9�Tit;Dw�ׄ�{U�9i,i�h�h�e&R �ʡp��m=!st^�9��m�7��{H�M�ט��j�R�[�S:��,G��Pf��ږ� :>��؍J��K�����o�b�O3����*���=��{It��<�,7 ��N���q%�5����bؕ��R�mqM��P艞{��
���uQs���g�:��|^ʕ*&�dN�#�_t���������
�}����W�b��Ӳ��.=�?��D��B�+F��2�c?���w�]{y��P��djEmZ�NՕ�O���'�9�*?N �گm32�J�<���C���(��1n��]�?%��:���KX�O���^_��.yкg}� Z*���ԩ�/���wS�*��&�uMW�-q;���*�$�쀤�{@�7rG�e�ΚV�V�����K�k�z*o'�y.�.ռj��HT����i�"[�b��N�ߊ�f{ssM���G>�"L&p�Z�/���:�B�*��4�R��J�Y���'��>�/�����ԋk�4�G���ጾ�� ���j�� 9K�^i֮aE���R��u�gaR�ۤ�.ٴX��[]6�Ъw�g7�{cx�~�`⛈4;1C���+�������4sn����O�:�����ն�]wI����ĝO�?%s�x��v�Z'n`8��j�R���5��K�3u;�-��NFV��ZZд�@1ǈ�ҫ�X�	���C^Z8�M,�\^�F��}�c%� 9¼ëR!��s�,2��n[W.�A�~;�8�n�Fh;P�5�bK�hE*e�[��7����{��2�XU��sN��.jv� ѡ�.�����Z>C�ĎgE[�Zҧjs�����!b���ڵ-I`s�wן��y�H��κhU��:��Z�g�cO����XDvXE�KJ��QQ�}U+�Sy~��!x��{f��k⽵���P<׷�r��9��AW�mz:�%�[�拨�n��V!�z�4��<=��R�ɹ��e�G����\��4�1�q]*�(ঃF_tDu={j�uB����=��GiϚ��a�=����}u�Wq��Р���$/g�=ܙ�O�U�f��^�c�w�j�Rѧ��z�sE�MA�5��6k�a6��ڨ���[`�uQ�C�6p>�b����� 䙉Q#��� ����o=�����y�;F�d����Mĭ�Vg� !���S�+3þ?41��6O7+��>�e��u<I
��e9�i	Б��*������f��o�:�e,>�P���PTk�r�F`G���qnYQ��S--3c��Xan'F��f�SfN#��~��Vfs��<5�����q�k��V6vVOeFg�X�l�i�����*����>i<H�^���i$f���H�I�ʣ�Z��4�ds@.�F��i���˒	�b�&���l��Q���nS�k���i@{��a̡L����mN�:q��W��;F��e;����~�{��P�z��%M������Ɍ�MĘ�����!��������6��i�z��T�Q�\
��W=�|x{�2K� T�:\�"0�� ���X`�)��v����І� ��.�Uk���0�����N�L;*u+�iQyns�.��V��	��q��F�����]���px&\�Ju�T.�s���k;퐻G� 1^�r�@^�r�.v�]V#(v�ѯT}���h���{Eh��#u]��R��ӷz������uT|�u�w��G/j����^�^��ȝ�m�guRލ��>��УZ� �F�3��{��%:�����R�Rܦ�oTV���mR7����t����2������Wm]ǾWl������V�C�y�B��G���.�I:jQ�.���8nSq�Nb@�tq�KN�i��\_�(�'�%����P�+x��·2�%[�:/�?��(�7�\]�N:|��k�d������z�6⽪��x�����P2���f!rݞ|���9{j8�"$�����k�Ot�gM7[uƙT�W��z��?YJ�G��<��0��a%
�m��ה!����5O���Q���vƋ6m Q̩N�q��8��&z�8h���=�O�.M3��Y�T��=YuZ��E�	��T�����)�;xR��Q��գ���~��-�K_$6F�%O �M�n�2B2;���~�7	�of��Z>0���O��#@�����v���,����jy,�n���f�<.qܡS@�B��g3��D*�򻣊�8����MvTj8�[��1A�x�W�Y��O!O �Zq(�:��l�����L��[�S�lۢ�=����\��#O0m�Z�߯9$� �C�5���Z}qD���`����s)��l��*	�f��p�� ��@z+�����zɏ��$7s
�c�%>�z[�Q�҃\�nx�[���=��@���2� �S�*�� ��vA�1��#Z=֠sj���g:z������_�&6�< �]���gF�e(��IT9���-3��SOմ��5
�z�G���!35Tn����eR���U��'d��nѹ|J��s��L����T�5��5R	��!v��7콽���M�R�s�q�� &L&U�����lW���.�l瑡<� [!yB�Y��i��,��!T��z�uM�I�<�#���� �#�P=���8g�Ӻ ��9��;��=Ԏ%jO�nip?�!�us1[Y�?����@q�m��c�o(��~�.� h��7M��\�F����[ٌB�ǽ�[]Z�u2���n� \xBǭ��s�� �x��,�W-�\�(h�r���)�#��W]�ifg%A��jC`̘ۂ�^��e̓;�*��i\6�Z����cl��8��ؗ�&�wu0�,F��*��T��U�w�M�:���{^��V�z"�I��� &�*L:5_�)5����vy0��qX�=o��X5�G�_Ӧ��﹮�u�t��m7��>�[V��eyZ�Z�������@X�G/�k�Nڻ�K3R�5-��f������*ޙ�gjɃJ���!�'�ʨ}ִП%���?�a!�*޾�錎��"&"w�X%�h�[��^�ڑ&�iV/:6\`i����K�*u	m{���1�s��W�p�;	���T,��v@��c��t?����įz�ڕ t?l�����p�J����\� N�~K��c��c�bB���<�\)�����_�+����լ�����;=�7a����I��KZO4.�e⮧�~���.�{��U^(<i��:+�G[�m=o+��CƧMՅVgkV�W8�/�⯮�ѷ9{Fp��U�+�ϣ���5�U5m)��o�pL:.�Pa��D������r;�xJ��2��$6H�;�(�Ew��\(Wk$���DpvC���a�M���gZΡF��W���`� Ȁ=bWM�I�X�>���R�Y����6��0;l���;O��>�Wv&��� =S�FSO.�A�(9�� �n0��Kg�\9��+���jx�m6xu�AA��H\T4g{��]Ox��]{E�s�ڌ�ׁ�N�SU�z-��w��N�&�.���ͬWt2�2v��M�U���*Ru*FI:�W��1�Y��RҰ9d�"
��f7x��S���0�[���N�9r�$������o��� Y#�5q�aE4�Py���~?r�֊P�<uW>�K��`Á�\�7YDL�9'V�Y�{�:j�Ӫ�hH�wZR�� x6	槑X���4�:;�/�a�m������W81��
��]Ӥs�d�~+m8���� 	P�4�9�t��� �e<����sW�E�/j��4�2��=�?}8������:C���*�_� @�� �іf.���aE��wt�>�f���#y���bo�K[�Ԏ{��{�k�NGjwoN� e���lj��ni5�k�8���(Ӊ�PsuG��H�Է�[j��hx�u!�6��+�����Q�����Ð?�,w ��	a���\�1£�Q��]��N����΂�8e����*e��9]=�\�I�=�~�]��եN�
Mp�I�����Luм/�}��>�_i�m�V�e���斷�yo���%^�WbU�H��]͉�?}��w�56��� ν|eP�g��<�=� ^�����;y�S3����E�;J�g%_��H`�*՝���tO�h�,=�nM�e�Y����j��[������H�Tc�k[�F_(Gs��e��fx.��A��Q�f/�����]��:L	
���amhȧA�|�ȶ�^*
T�r���!�'�����9���vޒ��[ҷ�F�2Ҡ�ƴp1���H��F�\ׇ�Z��D}ʷ�����Fצ�C�s���=eS��th�wh�d���'�?��8뙿�Lk�(N���o#i>���i$I�<a7�gц<�*5��2�m��G4���6����Y;O}�s���T�4���5C���]��q����~�Y^6���5���6�#S&�
jVW�D�	��Mwb�h�(�;]��TA(qCn�y(#q��`,�*Jv�*5x����I柞��l6�Qu������[�r�x��� �u2搲m<>�i�������P�U<��B�|[�B��8h�d���`8�YI�~Z�;����Z36�#LB�f�(Y�
|�F�����O%��,��_��PвN˲�
k'%�q]�H�2u8(4"��Y@��)N��(8��h�9���vE�j��|@<P�J`�փ�WM�_���}	�Cn�3<s�S�Y�;��z�(k��|�\:�39���B,�О>�Z�PO�T�y(%eQ
T�Ts*���
��GT�%O �P��f�Z�Py�h�<i(nz���9�:l��p<U��(ܦR��o�_�ۺcí��^�z�P�w���B�R�:�ۇ��)��T�6TX�x'���.t��%Q���=���Sc�<6�N>j�YE�=����Q����;-��(��vc@땪�e@ꐧ��B��
y����
O%�5��DB���#������%7n�%�վ�|P|T���b1ڎq��n�� �-Tx��U:��=�Nh�2�����Kp*��%2���XI5i�u4�qN�]�*-.�2w)�q�)����!�����쬠5/���晅���JA�q�m��G J�v���T���*3|�����h�����du��k�A�u:cE��j�wP:�J�G���!O �Q�A�ҧ��5��S�Ƒ�[�@�5g�X�(멣�Y默
�T�: �-�@_����+�b�n[̆LlB����}���mp�}݁�q	�����7p�ThT�I�A�~��=��y�6�C?ۛ�Xe:��O<N����֫+W'fi9�i�t
�ޅ�G3<�p>�pz!������ Ϣ��:����;���]�c�
5�`�������<w���T�@�䁑*Bג����Ӊn�O���j�B�`)Z�F�D�)�[%<fDG�g�<Ui�}g��@�D�{V�,LU�u�:u�Aڦ8��T�\��J������o��/������	����t�M�� �5�\�ĎB���}Oh�pE6�v�1�T� x�yjNh�U�2��i��*��ˇ�a����� *Af��}�Vx�nc�3#��2ڮr)3L�Ͷ� ��R�VG�^P.�`=ڤw�R����f��t��XV"�{F^��~h�$4��D)����B�{�B�y��;'�<��p�L&5���B�2�'~: ���m7:?��*b�3��Dk�!*Q�]�S�i�tʙ��T$n�.�kk�.p|�;mK�2�PpP�%v�;6<�rz���O�-#q�)	�㲩�;]�[�&#����
��;�ŚC�R��z��O������U6�u�gi��9�K���}\��:��]�{|�ԋL���a�5��fJr�<���x��˂�uT_1�{�u=Ky�W7�����'YX��#Z�;p`V`�U�[�۱��*���ەŁ���VZ�&���io��W��0�A�^�����!�C���[�g��%߭7�b��2����Ӕ��.;,:¥Ӄ�K3��|U��vR��~э���S����r��m��L��fz��]��NK��Ф���<@�శ5�DwF�5nƽ�e!�{�`��J�-�Tt��t[+�Q� 1�������h�E��}�s��1=d�0�f{G���u�ڙ��sL��A���9�x&�q�#��A�9�P��Lw����UVj��R N˵q��>h��G�mG��x"��L���b#�4T�䟫~�/|s�Ä��Q�&h��F�ʧ"�X������Od\H
|P2:�����;�ǒ���A	�ΣN�JM���Y���>�d4e�Uo���웧�uڀ�s4�r�Z��׻(!��������-�uM}�VZ�fY�32�nk6Gf��'��*�f����;�T}Q��;}3�^V���u��s��Z]}C{���z�,f���ץQ�̚8Ƀ�t�Fҝ�_p��뺭���4�9�]}}��~����Ç�T�Ve0^ָ����_%�V}zt��Z�4�@�a/}*y^��#�9W؁� )�vps~k
�(�:�?p�|yf1�*���v�-qݺ��b�m[�w�	o|�����(�����}J.�E�cZc�a*a����J�-�ҵҀ���T���\��%3al9���_S��e(9H���ZѷutL@�U��I��I�o�B^�9H�'ӥS.\�ӡ��ɐi7o׊���4��C}����s��>�57U.�U4qgu@����6"t��������ˮ��˫*n�!�ۛ�b��Uon+��v�������y�v!yg1��Dʷ!��sa���Ԁ6�Z����#�To���8 #oUV���|:�t�v�o�!��Nc�U��������=6T�o� ��}Ъ�]��麩p:�0 w*֥qH�i`�uwJ�{^�.�C��qrꮯ��0&?$1���O�Q�[���-���3.1������w(�����҃pH�G?�6�Vi�F��{Wi��
��l�\\F�M�n蹯���B��vz���1���}{oݥR>	���V�C�4OѠ��r���9��c���x�ڻs�T��b3��5����H��l�rT$��Z�L��G����#qP��<�U0�S� �<��u���TNW*�d�U�?�Yi~��*ޔ�����9�pX���xi�L����Y����*5����3?%!I��2�q��p r�J�Ѷ�m,ť��յ�oj�;]�Е��up����}�Օ�����H��W8eKK��g�� ��5�\Ҵ:���F����·9����kLh>U��{��`�)�H}Y���\�֙�ڭ�69H��M�ӣ\�0�YӥU�3S�r��U�4���W�������m��ק���~�i��q!\�w�R�mj$A,iǊ��}�
�bi���6���:gs
��ֵ{2L�Cyk̩
y�>
Q3
t#�	��nc�8vc�w]�F��[R�u�j���
��?�V~}a�H)�q�T�K���":��hB��O�����:�)<��q@���xf��"2��pXSrb���s�N�}B�֭w۔��얕o=ڎ�m����V$������nk�Ѩ��k ����ƥ�{��Q�c]���5�\��k�\���	.����ՍՕ�mN��0g+O����v~�T��C��
���1{6���pi>?�cj2�m�]M�hѮ-��e��u�+�z�X�×6�t�U��k�0l3�NZ��VC-�����"V:I�� �O�B��*V�gm:/U�I�Q�v���T�/.��T��>����V�}\Ǐ�� 8�]3�"5+A�"�I�[�e�O��G]4V�?�=5�t���-3�px�Xk�+��0G/E����}Ep�yk+�J�zV�4��p��� r�a��%���b6�N��Wߢ@3���Xvu�W=�`m���{��*���n�V�sZZ��v���*լ���o�$��L��-8qXAN検��)�MC���H��,_�6�ՙ��]� A[�vmV�ÇkY��|r�{U7��vY�U�qF�WT��1��p>���,^�k�T{܌I�R�Q�u���:�)��N%�:��T�b�!�����lT�*'V�a��y#�SFQ���A�D�TuHS�j�Bs��=��ܠ �Y�9�ď�I'���y$��E�*{�q#��>�Χh�ռy/k� ��<��D}�U{}ڎa��R�Z�v�*����0����s,�ہ��J���E*�k$���U.j׃V��Fٿ  @���������	�n^�Ws�>+m:�j��@Z�U<����)@4�E�?x�1柘;T� x��x&;E@�-tMգ�N���>���7�ג�����e>(S�O ��ak+��ϊ�(S�`�|�'��1���e�����ƨh$��<��SNT�\�5<�m<�2�SjJ5@q����aL}���"� ?@���h������3G5�Z���������K���$�e�x���×��4�Z�	�Js������l�����f惙���� d�.w)��2�9���uO le2cTTx��D�Lu�2�x�k2a�Q�������53	����s�pU0�I�2��C�v Ǌ�iuD:io/�n~WIjmM��O��3���Z �7���LJ� k]�N�	#u ���^�\���s����k��gY>
�
ڭ��$�~���H]�W�K|�8�ɳ*���@�����O뚩�X��o`;A��?� g��d���2��s0i0�6:�˘TL=8ju�8x��HM ~�i9F��'���ޠ8�S7����MxuITiS}P��s<�[�4;�6-l�	��r̹C@����Z�og�=䇺F�<>�SN�ѦH�ȃ�7�?讃�S=��v���O|�-�*Bג����YZ�M����s!��<U�����9�>j��7��s�i����^�R�ؽ�-c���Um
��f�]���a����"A�i���f��6j�q?9J��B|�i��X= �]�/y��yw���A�;*R����6d��p�I���4s2���UR���M�M�y���<���HV��ڮ ���#���R����: =�_�-m<�h�ӎ�yB������ Z,Z��ʠCr5�'�i�a�s<z����!>C�yl�5���k�5����:+� p��X�n��#�cv���P�ȫ���"ʍ�D����|�F�Yz�����s�vʔ��4if��2A?sO5�� ��ٴ:k��r�]��[;���]�'�C� ��1R��أ�B������eK�'�S?iZ�� ۱�ddj�� e��lg���Ñ�~�P��v�-Z᯴�O��>�jcͻj�ޙ�����!G�x��5�yqTΉڂB�*p\Á�s��Z�9Z�� ��i�Q�S%ü׃��*4��t�*�4[�$�3�yy.�4]U�/���!��P���(�E�z�1'x�Vr��~j�;6o�p�L�Q��. ��cUk���kHI͘L+Ƕ�+��f����9�����͐�Q�����T)�G[3��+w��ү�����L�:�"�:M&��a���hW���9�6�u�'��x˔
�j>)�5YurX2�Aׂԅ�jvMͧx��f&U��k�-7N�&xl<�*����7��ZL�Ry-Tu�A���(<Jʢ��1k���֤ESަ$p�ձ5nQ���|F��O�n����T.�sU��jK9�$�
ɭJs�&�Aԅ�h�&�+#V�O��G�dN^'��X�m�w�}�$��vO��}!L9�]'�?B�ޛX$�`�+ʔ\;:f�;h��0P�,s]�c�J��w�V�=��U/,�\^w����݁��-��sU_LQ�2w��<}h{�u�
ܜ���SYTSA��q��V������X����ͺ��:fz��F4:#1�ɢFm�`��'�M��U�9�纎�
|�/�ʟ�RWi q+>c.�T��]U���	��3��۲ܙ�o��ѹ�i��p܍��0w�)��D��R�k �+;����wV�'ߍN�q�F�x����uy!���p�?^K�/]����ˁ���U�]�{B�~I��}�� W���tr���n�pب�USWO��:�ɣ;c�Li4Y����h�U�vR�4�>��+?�:��S5j���$ZsO���:<���G2�4x��5�D���4j�H�w�!�l��]�!���>|�p�Q�&<ѩ����/hY�l�ʖ���Y�5�w��(=�d^�h]��8��!RJ����$+Ffr�i �*�^���Ъ��L��K|����7A��-��B�����P�U*T����Pg5
xG^B�s)�F�z�('�@�gU+U�}�*Ҡi$�<g'��ϝ���g �p�G5F���_������>�(8�HRy(<J�eR���ĭVV�`�Q̠ޣ����-V^j��Q��<���9�4YJ�8��
O �5Mc���VAĮ�^Rz����D��y,��- x��9�TJk^l�S�:��D)K�Xk}�v��Ũ�QYg�H	���x�+5n�#�>�״n�w����9��8���v���>���^	�T�'�3����L}�������D'�Nsˡ��,���j��+/���x�${�Z�躧
��<�=��ܴ����k��w�sA��4R��q�x5��J�e���N�����Y{�&9-�����(���*y'��w*��ف�]�o��5�V�9�"B�Ox��*@�S�?B�>֓N��9���tڴ��z����@�*�ޓ�8S]��+�.�0�Tp��ۓ��X�$�ձJD�}i���&7��3�F
v1|��e� w�_�/�._<5L�����O�_��~���p̰Z�ژ��NR���Q�J�X�����ٚ$�Ѣ�.�jys�wn�4�9a]Zb��R�B�PeW�Ǩ�=�m5�eS�8�;�kF���l[��P��'t�$MG7��_�8���{D�:������Z�q���W���2��k�+���?W�7ƞl��ܛ��C,�Ǚ�/�F7�̕�Y�Oy�M4;�������y�}/�h�j�=1�']������{�~_�Dޛ޻\��G俍1�����n���2�������_�7�0CL�U.�bw�L�����%p�D�w��j�3hx���()���:�4��B��Fl�&�L��ܾ�ZY@����˻��{� ~K���3X�m���/�*���<�M�d7'ÒoK��9*]5�1ِ?%�OwY�4霞J���ss[��-T,�V'gj��7(��ĬG	���Б�����T�fA�����:�B�F��ɕ��j!��y�O��|�Q�'Ot+���W��ę r�u���K$���\�5��FW��M��ny.�L�$l�	u�3jC�*.k�y��r�j��j�{���+D}꥝:����q�����U~�P�9>i�
q�Ϋfw3���j��/��9��+�8�H r�N�C�O�uwQ ;��!ܓ����{� ��U�3y�fg? � �S3�^	��@$�-4G�&{�Jv}�_���Z� �X�]�V���5�[SkK�3�*64X�q#��9� 5��:�0���t���׊�q����}
���b��®n$��	��Q�Q��2|Sp����2����F/_��D��Mg7*�	������zZ5�|����B��Z���8�+�E})N^���I��	��[�V9�
�pu?YfuY@Y��G2�#N]3#�t��b�cC�ƻ*���x��8��u�U(��wB��漟��Ϭ���@&x��VC��9��N�� ߯3ƍ��وh�y�%08Nh2�7|���6�t��{,��*Oـ"�4do�!N�ـ)M�t)�7(	�.t� HS�������ذ��Ż�w۵�A�T)���ӹt�+�Ԟ�jZ*6ti�gDG2g2�.�  �̤��f��P�{��;�)���殙>�S��
��)%G�%�X����Z5�D����zOާ�X ���\�KE9����P$l���IY }�b8��r�Ĭ��:��,��	͖������ #����/+k2㿚*�1�T_��U�h����>*\x��U`�ϗ�ׂ�G�3N���)�(��:L�� ��(e��x̌�@P:ʨ7� ���Q����1M�ˣ��O4OH����#��2�����#7�����1� �]�#�u����܏�{�x5�|&&걈�]z�{����a�,���GPpu�)��Ԩ(����&�-&^���0)��u\� 4���-��8�70��絮�ƩÏQ֙<B�2�F����g�h�B�R�"NC�t�T�˶���0���qf��I�SL��6�1O��Cn���z�ͤqX�9R֥J^x���Pl�O� Ҭ)M�)$w�O��n�r:�dB�q�*yA#�k�R� &������k\84}ʠWTC�����ݗR�U:��r���e#��#�:u}�9���p��3����I"5N 	 ~+UM��n �]� ٶ=U4��b4`O��k+}љ���p�y�A���%>�Ni��9ni��B� ZS�!�4)�:�;�T��X!��oeH�ﲮ�
{L����GqZ��M�?[*����F�h��C�����w�6�R��6j}���G�ǁh��������=/�C��pYHS-Tξi���@�u;�%L���d���G�q��\!t�=;�#��9��'��UF5��dm�������+Gf�H�`GV��ۭ���P����R?RƓ��9���UJ�`h������EJ���+f�(�DB;ه5��Z_%X7.W0:Q¬�E�w��g2h��B8e��v�&��w�����Тe�Y#T���eU�D���lW�s� UaL��Ln�N�\vG0�_a�+fp�P�͹�f�=�ZuhT�=F�X�i��oI�`� �)
O$᪃˫^
�'�]��O�#�Y�v�T��6�&��5gG�����@�^��CvUlA<��oL�$�0��Ytj8�:�cE٦[
��O��ǇLK�#�%9�e�VH�ldt���5��L2����1�A�"%�TBa��?G�qY �ފ�FӒ�b$�}�~�Bkw��b�qr��g�]�9!Na��u#�j��r�I��ke��������A�={�;z��/�>>~������gc�W�_�?�6�i��.�	�evX��P�?r4�gr F�����ǚe�(>�.q��u�!���}���5c���u����k�=�\�ǒ67����	�B��ԝ�mAUi\�i/iUz�Z��v����uAH�Ī�T���x�^�p�n�8�ϒ�Y�*z��Y�5
@�jq&�e�g�P"<��ދ2�h��L��V5�nx,:��S�}6:�� �p��9fA �+�ݢO�A���M���%EF��j�����n�%��_�;}��H�_M�p �˂��f��m����庌���D癆��%S�v4��
���{���LɢZ<GquB�AsKu�	՜N�B;�!t*ڙ�闷1ϧ�h��S��������9��$+�Cl��i��r������1�"�*Upʭ����w�[��Q�o[0c� t�U�K+�{��ͶX	�6fy���P�4���;Y�����
�A�I�~�g�&��S��$v�YF���S�;�h�hX�&�A��6�+�,��ZѢ�.)^�#��.��t��GqIõy:��X)�mn��G4%J��|tR�%�3dc��<���ZL�ʀ������\
{���wEf��`%S���/i��yKU>�Yi�ޏ�'`8Y�ִ\Cc���_�?��n'-���pl�Fp�j��0�eLG:�����miϗ�U�7���uJ��y�?%ui����(7<����Uð������%�Ƴ���>?����z�e"y��� %G��I �|q�������*�i:�2~�$�.��8vU��!���.�z|�ĎG�v�Ч9�E�At���h�lJ��׹sF�N���1��{�۸���//N���K�ϊ5j���5kZ����vod,+��i�k.�\�������[�n�R�`����a�B� �#ER��Plp���M��cY�L�R�X�9�-C.c^7�B��l��vY�����n�y���ȏ5�Ǘ��3�n�4D=m��A�T�w�M'e���eV�������<�2�c�]q�\r���H 8F�v%�6�u���M��)�ә�T�Eդ�k;+��׹���3�OEqoe�b� 1$�+��U��A�t�� /���Wy���w�c�t�������:]V�@����=B�����J/c���].�*`WT���O�����6#�	��+��`��U�e9:��tˤĮ�oJ�ѤKA���|Ph�:�E��y �&1�p�r����_���z�3*:���3���ӊ��]F�c�rh)5����5���S�Wv�Ƣd� �ު� +|� ���͎Ԧ����LH>\@��K�nh��+3G�Q�U
S���8L��P�B��j�e�"y*�.�C������O�����D�E��T�OPka<�s�?��Ǯ�~�J ��{����̕{�T��\\I'��s�����IOh���p+�"��]�q�\Ff�?�\2��p��)k�������t�z�-$���,L[tD9�*j�ؒ�ῢ/�q^���D��؎��f<��ʅsM���8zXUǵYѬ8���$=6X5GT�A���B����C��� �k�F�b�+T0K5:�_����b$���]$ğ��&�_��L��++B���T���d�D4���/�Y��g*IX��)����bm���_�ʭn'_�R���������@4�Z��Ae:��1�#�eoQ�Y�j
�Z��;�Z���
�+���gA=��+��*�:�]�gv<N���)�"g��$y�rA��L�Fа�S���{j�.,ljO��A�P���$nJ�Q�5�A�^e�m?�c�:�vT�:���jx���6���Xy�J�AUZZ���}N����m,Y��7](�;JumH:�\�#�X��"�~�3�$�!tƠ��m�_�N�ec�k{�t����ǼЩ�$n��wrĝԀ�Q̢˳�2���Z��Vf��*y'o�5�+��/�k�>�Gy�7�8��*����Ж:����W���8(����3���8i�,7�}E������=��$8h$s�7.�l�8˘aph<��s���)��iR���-��	X��Q� �y���F�cVy*��k�`�f��&&�a�vUZEG����{�_4��?�p�� e1�@���#����7���+S�:��J�FbjS$�V���*�zx+�������8�i3�3�,V��l.��$�vV���n�p�N�ަq�Vxd�y��Q�W���gMӗ�����syM�����lp�yЖ	��AЍ_��%7.���Ȏ�����g��
��(N���Y��Q��߲[V�ʛ��t��u�^�߾F��.+�ocG��/���_x�V���&Ӧ�c �"b6�[�oV�x�{��������S���@�Ni�
�U�"�f�s0��3B�	q��f��t� ���S(k�T��L�k��4�`�N��"��vnd��<%���Z�}>�=?��bZ�4���D:v*9�!9�/+&V�V��.ܛ� ge�a�m��Sp��;,>�eHcuL9�GV�r�̂�M���gAkߡ;벭���'�t��e���赹�5��S���:�y�;,�i���"�2�e�H�L��0S�-Ө�"s��ɎHz��u��h���s�̦hc��N2~�oy9�%w��c�}����[�70�Z�d���j�{�x��ܮ�~̯0l^��wwXC�t䥮ihn\�|
��5��8{Kze�$����F�Z5�F� µOh����q@��鑣�>k��}Ju�r���u�*��?u!;��Prėl��8����e�DA#���N���t*����a�ft�7��n�\a����EݍWK���||�������5�p9Gv׫�S���'�����V�͝��Eko.g-4�wZ�A���0ؒ�QiOy�_�*b�/Z�Tq�ԣ��y�>k��Gu� #��}T�7(0<>���8�Y� ���Ѱ��<��&��$Ϣ��M:��Ӛ����;[�8+vѽ{Ǻ�o�И}V`��p!_6�k�㎅t�	e�*�k'��
�����e�U:�Y�k/ ��%>
	��']]R`c�.�6��qU0a�tb��nAقtU�v��e��X��9��5p��uj��*�LeV��.�&a״E+��b��j�:x�]&蕽*��unZu��7� �z��74	�ghk���(�T��Ut�Iܻ�+ ���7V�:E.՝����P��Z��snܢ =����ᴪ��;1���n=��/�4ss������i����&�F�����*}'�(��x�q�JwJp'S����-2���S��n��vzOs��Jp��������2к^�ڙ{s$����&�1���Q���Nm�7�f��Tڍv�|vWT��T��<UJm#!� ��.�tJ��M[a�!^��m�料G��o4[Va�%a�����=�5��5�JeԮƹ�K���w��z���\V�;�o>���t ��T�E:�d�G�p�uT�ԙ^�q�\U�	;!U����qY��Y�̡Z����jtB�ڽG2�j͒�v�iQ���y�3	���{� �k��rI]�O�wĮ����	����1�Cx����F�����/,����cxBf?z��p� �އH�C꫼�����Lj�i��'^�:!���˜���q������:q��z����ӌZ�-�\֝!�{�]�����^�U��~)�u�0y����H���ԝވ�O޿��֎\�
릸��[Z�.����A� ��g��?��;�UG^~� 6� SRW����r@So�$�={�TT0�$3��9� ��� �� �� �� b 			  !1A"2Qaq#B���� 03Rrs��$4b�����%5@CS�����&6Pcdt���DTUe���E`uVf����  ?� �2����� �Td¾���?]0<I���c&��O�����2aY1�zD~�g.�3a�T|Cި��}Pn���}��N���>%�D|S������/�#�����o}X�=�c��Վ���#G~�t���{�GE�=�Y����3��t��5}C%�C5}C5�C5}C5}EGƫ���}EA��� 0���&>;�c�O�1���1�ޣ����G���~�A���T~�\~��"?O�?	@��Q}J�_�8��ڏ��ry��
٘[����W?,@��V��8�r��ee��G朶�^]o�0�rQ|#�%�0��5h������;�0˥c<O�{w��J���2%�^e�q�n������j��^��[�L��n$�o+%��R
��Õ/��W*w� yW�/��K���z��z��-W���y��5N��>�=ZFuꙿQ�������?��c.�}��GR�M����q���8�/�O�4m͠�qϕ+��_��t<�YvŽߩ�2aV�*�p�9we����X��ER����c�z���tgꅗ6����_����į�5Z��'��RJu�x�{�+�d{�g�#� �5����վ��m%G/��ז������� =�������� 7_\g�u���r��z���h�?]�O���|�R?S׬0�v�u�p�W��1��9uta��*�yU<�]g�x��Eh*@Ęο?����� (*]'�X� 8����� &pm�s�����������4����2�L����u���>ȿ�s�z4��ǻ���᷇�� v�Rz�S�Z1���Hך��3�I�=����Tb]h���i�n�Y�E+��1�M!����h�����i�F)�7�BM��(zð'?TrYٔ2����}���]�����n�h��?0���¶�������� �_�)2�$-��ʼ5D�4q��f�U�Rr׶�����<��	f�.��Ԕ��K�/�nvt"��bY�i�:�ψ�|^Vi�N�B�1�:òU�V���C�!3�[���9�����K���g���|���Hy�]*ї�iA�e�vڛ���y���
�t���M�H�䰙��7R�Q�*7=���Uk�34ey; �V�.��%�V�T��(�.�w���tj/�J�J��=�EӘ�`�0s�E����tT��-�Be2ԴL�)*ܡj�4�=O��O˺��Ɠo\c.s ���Y������!���d$�jz]�{�0��&m�|���Y���n~m�&���A�-�e*�J��eci��m#���x7��n}��*��^��M�QHqĶ�%�r�<�-�,�6N�#�����㘥M��6{���施��֕�¢�;��8��Hƾ�ů'z�YQ�Ū��i̸��(JuQ&�M�I��;#E�%��\��:BX��fU�)m�% ��3ZS�aK��N�}�d���;��Pu
࠱c����T�"eg�ڵ������<cg���H���F~��_�$ϒ�2�����>�*����Ŝ�Kn�/s䶋��f�m�w��Z�
c*q��I>pu��krI��Ҫ)AW�FY�v�ZHMRLx��L�<Ooʉĥ���!*��t��"�n��]Q�]n�p%�(w�-	'��� 	�.Zha��p��ws���� 4�.� �"��@�T�e�����%*N��>��F\b�^����Eu)t>%2���!	W6�s��&��0��$�Ԕ%-4����0��j����uL��T�U�Y>Bcx�v<�Iy7�_��Xnb禅�Tn/R��X90�[NJ�AI�_�H�3=8Yf]�ed��<��qdf���!�+Prwtԣ������g8��6��@Q�e�1MԦ,�WAĩj�JR	�C��m˷��Ҧ�\�09���'%a�W�ĥJy�i��2Y�deZm+Km�<�� (�'X��]SMV�)qSrHZ�-ή�*��$d��8�jX��eX(���U�I�HJ�sG!�eg嘜��8�t�t�Ru)QB%�����~N���6BW`�{v�%a��I������(X�&'�{��C~�[�PChp	Bt���ag��e~�+rd����G����NZ�R]VG�#��ʹ)q���V�0�W���J�t13A�������q*뽴�=���;F��c�Y�>)�:u��L}�����;1*ۀqi����쀔�ciJ�,�  ����9�ܑ���B��b��s��1&���.ʬ�?��̘o
�t�����jjS���N��>C�3��*�g�?�P��6RLL�۞�nNqgx����?d52���J4s��m"�Va�l�;'���*�)��2�5�R[R�Ad}�NSܠ�3��]I�U�n���#/@�t��KJi	�H-��M�<cvQ6��&�ԕ'9����/r��D�[(��lܰ�	f�S_%H��Q���ק��S��<C
���M���oS�6>����S�7$�SeC����쉖�j��9K	�g�*��B���x��jU]�����
�.���{GRmμ��̫jęvS�qe��a�R�U)���Ku�%��7�8�T�Z�/�:�fms)�Y��r����r�������f���ZV�l��H�EOe��rO�t�l[d��G�L'���&�>��@W�)(	f��;2�f\�\HQZ'�o&-��'O�0�6�,��W��b��W�ȟ�u�'d|s�Jy�Z��S�R�+�O']�7h���3R���z�cq)ě���&>�^�؂��������<5o$X���u+�B���v(ײ6�u��0?���D<o�?r�}QN����5o�a� T0��#?$� `����M1���:�IA}�6��JM��N/�%%cB8wEbV��t�r��۔i��T�Kd��-~��MHޠ���7c�oRⱆ����-�.�X8������AI�M��_� �ey^ֹ�%�j�����G5�n93�|Q����ӳ3����qjq�M�|R�ǥ�'-!���`�Ʌ�ˡm���^ѻ]�7���
u��BR�,@��qꍌ��7(h��w�T�{���E�����&$�Ҫ"�l"aO�>��دw�|��$��gev�Au��:ᄿ$��s$���<Dm�����^LM-�L����mD @M�]P�l`��.aW�l(���t~�>1����d��y�$]s�X�q@��|���7\Lp�:�a���XB{p���y��c���7�I6��:�C�Z����LS�r����/{)I��`Q�n�R�{��0��*�H굷baٷrfU�_qG$�- �3�ξ�T�\G�%[���_��e�djt�ۖJ�m�_�.p��8�335�.㍣�II�b^��jx �!���*�J8
Ozx�ɥ�'*��ۨjaK�J8�w8�|᱕��<;�����(�:��r�P��r����*/�-�tK4-d��y(�/����	Զ�/>�Psr5S���	�@��)��~*Ff.].!i�n�HR����fRD�n�Zg7��K�2�Ni�.��C��ڣ���aD�V����hз�=1/����R��M�Z�dhU�7�+x���:ҏŬ����t��ܫ
���x����z�ja!�*���	�Mj�u�l�����-�JN �Z����֒!�r{��q�="�G0�(S\�DK�4<l���8���n%\�@����Cf� 1.��R�m{uv�,����:��S�BVc����B���}���*)��?=7���R��D��[���M�Z�T��r��gtk�
��@��|�d��1�.��o� n�u7��0�e�q'�l})䮵ZN��� ��°�V�ʹ6�� �	GP���;X��aUF��НRF�)�J@V�xZ�TUNIL=6YL��i)�nը�&�J��ge��LӁ�8���n/�k�*�G�%��>U6��v˳�@���0\V6r�Am�jzݓf`I�%�6,wkm7�IP��t��\��d�SO
+<y��q��=�od��6$Щ�e$�i����J���ck��5֩�!�&[*�}�]�4��J3 ��Zv�J�n�#(�:�*mM�(�O�O4KUߢ38�SHm�N���)6$�D��g�QM}հ^CCvm� �V�`H��T�J�S���Q-O 8���������:��zOT��JL=7�cr�@J�.�Ll��z��ٚ�lr���(uKq ����@����2�Ίzݝ�e�r��V�d7�8��dy�r�A�y+p�]�%(�w	��f]n��:���k�P��������]��O>��d'RTt���//+9%�X��� vfTOE��U�s��h6%t9iY�r���A�q��zӉ��=b�U�'��J[Ϸ!.��|�#�u�:D&���츽o)��RX*�毢z�k�*Ztw?<L��n鵫J�����S�(��:�l)�����3(�����!"▬�:���=Ӭ�{2>)�!��:�f�<���iN�K!#�.�6��p�+e�%-��t���g���{��Zo4z�)PZ�e�I�I<�)�I�nYP����C|�6����T�f���8���o(8���jS򒌠\��Гn�{����O����kI��"YQc�O�f9P�Yq��QR��oa{�H�����Y�O�wY�M>e��XRՀ>Ӻ�^%h,UEBrr���8
��Z���l�geܔ�eR�%n���BH_�]���Ȯz�LK�n] �T�Ϧ8w�zuST�:g)��fa�.���Wc�Y�(oM<��V��q�pKx�|��u�d�r� ��^��|�)$���F�N�,��.K���m
R���'��[�)f�6�Ԕ�$�|�RY��;4��_KiX�t�(�=QZ�M.Y`("�
r��戞�lT�T��R���'�˙�,�Z�}�h�4٩E���Jĕ6�bcf�f�<��p4W�mh�	<0�zڥw�*2�e('v�).�b�6�q�$�̔����h]*IH�մrc����m����_�q'
��Rh�EE��C��5d8��.' �kM��A^h����9?A�̱/�)C�RqaN@���mR]�d���2�5/���1'�"!��m�~`�6�#
���q�9RC�V��兼Z�b8B|:�5�k�jt���-�6�lR���d1��^��n^��Jt���L�>e������>c�]A=���!ɪ�A��N�-%՟��M��%���6�ҹ�'�N�z�flk>� 4Ä���&~�^Ƞ�[��=��AQ��g�t�G6�P�xO%v��-�'V��RV^��H��e����}-��W��O�l�RH|1����N�>����`ﰄ�T��*',rn�_݋�J�߬�?ǒ���vʼ-�Dx�I�|�wG��̕�P�V?�ŗ-2ڭ��p͋�I�:�~�~	7���Տ�&� �<O�G9��u�K��j#)y�v�?���So&�ݗ���:R�TY��0��C�f�[K�Z{��q���L��%ٍ��C�hL��r�/,���V�N	MǲY�ڂ�wIL�S��a�%\�
���ԝ�)�Rq��i�D������+K�~1�{[ARL�F7�R��Z�V�ki�O��~J����~P�9����8R�E�J��(�t���R�0�n ��b������GW�t�r�E��%0�1n�p;ԕ�C�OY����͕���ʄ1H�M3,�AnY�\Bm�M�d'i���d7�K���\[���`��e+K�7*g�1kn�y���L>��hT�o����J�2�@��[�'@��"�D�u����>�.:�%H��������s�{K̦�P:���)/�r�ʋ��-wHuZ������=�.oL���c���Ҏ�������L<t�t�t�=�<j{�:���'��)9����)O�*uX})�BR�<G�[I��y�M�tK��Pn�\��J��J9��Z�g�		)JF�_������E�o�+�L�
��7P��a�%dy�y��RغՇ6���~�ӥ�$�6䫳NK7��k����k\X֫���%)n����];L�9\�W���m�W�2����\m�Zߒ���̄��о�'4��/����p��K/��yE��x���^� �:���K��=".�Ii>��P���,�����F�. #��1��lmy�����7q�\�7���W�;Cؘ2c-��S�`�Zݖ��-��	A̧p���Lˎ��#
���������}���KR�� wh{�1�Cd�c��}�N��Q�G9�M��I��k�ŧ샻CC��'?T|[9����:��Zb�,_�Q�F���L_w/�G�-f�NQ� �v��t'N�݋u6̹���tn�@Fig��S-k2 �7)�f3��?�G��^v�\JIwn���k�>��_���ŽΧ� W����q�j��>��RM�������RO ֽ����G��F׃D_��e�����4�2u����� [��	��#�� L_�J_�T_���[�Iw`�B�t���[_ډ�{��1/;&�WBe��)N���g(�У�R�g���i.�>b�q��z�0��D�o�k�5� EUU��-;>�lK��Z=���%{"�bm�J��J�#�.t���?���m|ƾ�X��k��ׁ�
d����J+�]�����%EK��}��d���TK}5���F�����Oo����#O��4><:F���?
~p��6�/މ_7�ȑ����g_��f~�Q_̃�:�5Q#������lK��7������36�`@�| <�=g���(���(��3��_�#��i~�6��;GG�э=�H�>p��Wr˹���o{�1��c�3�F+���'����Z�̞�7Wh��O���ӌh�ۈ1�V$�A�A�=q�_�mqm;c|���J �&�F4g|�g�/�q�g�I�&)T����o0���ƣ�H��3-.]捜iԔ�=�61�{�-D�rEI*!�n�x�z��E»5h������	-P*��$J��z� �h�g�����)�1�g���w�`a���W��ߥ6�0�����n���ײ3���� �s��NM��](�mM�C�@�����\d\�ۿv�)dty���c�3�j��^���"��JI��qC��g��O�A��&_y��$�dr��zR�	��B��&��%�H���1�Z_(~t���-/��6�yt��2����n�>N#kvF�Q:a���}-�K�%�l��8�p�VH�"�D�2�M֥��W�d�!���-*�y�a=�q��3෼��v�ĭM����ܦ�8�	$��p���jXj�������K[�[��A��ߌL�6q�UV��$��l��uM�1R����t��)I�zY)[u�ڃj9d�VP�b��g�;=4�?D���� �DvEj�ݒn�g�x0�ˏ6ˡJ�$����J\�V���r��ۖ��BBגT��rϮ*Δ�J]�����4�&���:�RuN'R����h�
 K[��q��� 5��ZWf(�l�㍶����e���R@D�F�B�;NrnZVern�u�2�I�[�P��u��N��lL6�� $�X�mm8Fx������/���>>&(����1��%{#h��+��ED���h�1�h뭼&;<�I]��9�x��m�n�3(�k�+���C4���S���p�[v��	:Z�y5"TnIFA⎫y1/:eKt��d�u�	 B���枦�Rf��gk�VBR�4��<|P��Bw'�a����~�w��NBpwww�$���݂������lUW���V�Tϯ�w������9�@:}�W�Iᅃ_�vw�(�K�6�\Z��������&���S?�K��c���t� y<Y�������'�Ӊw��r��N��bb�m�����;����4��iTfV����%�����1[�s�w2�È��]��T6sJ��v��C��^�W^����Nb3�	8St�<�SA������:7��U�l��+����_�D�ٹޮDZ<o�`���]ڡ�$7	�*��$p�5Ap���<�՞F�i��N%>Q[�!D�jf3_�l\?#�ǴɌ)7HO��G9<����_=��sݛ�R���\�0i<��d֠����~�%B4a�6fdm�tN�9��L��C����8��]�ͪ�7���ӕdČ�oel��5}HY�����N�|��{S�3�YV�x�|!
wA�J(�*n�Y������zE]!����)3W i�EG��*ΣW9������_���ݠ$���>i�tg�L*L�����L�[��⺰&#ٔ��4F5�ŉ�j��л�F��)����-s$�����'<Җ�z�W2%���1Y���E�V�G�>Y�?� �S
Y^:�>�y:�Ǖ~��6AH΃kE�����������F�v��v�cÝ��48��h3%��1��b����\�����[���;�[�Q��Q8ٝ5�_k��������Ƴ��0X���V����Z��=�ʎc���:N.4�� �u��+����a,u�2��'/�d�++##Xq�����!)I�� ����+b���Lo�f�d�T��Pn�16A�ά�"m|��;�!���
�t�����m<���i�����}Y�����eu|�Ǫ�6n&���K�0.�6~�cb�X5Q�{��lVJ�����_��Y6ѕ��%��(���.�p���cZ:�%j�~{�k�}	��-�D��_T���p��^AȨW��R$VN)��*o��(���a㧲��o��/D�ЗO)��V�A5���҉��M�%��6;/���ǐ������Z��ob���ru� ^F��I�Q��)����zW #��r�U$�x�Y��%��o����ъ��o���.c6�9j��?uh.�C�|�}�x�e�Яc��^Ʒ
i�Sfd6滆�L-�]?�>�O��W4��JU2,�T��3���C���=�[�,o���'*m�;�."yn�3M	1�ͭEn�P� U�������v�8�2���"Gϑv���a`'ϕ�[Vz��?`��D��x�mm���)%Y�����k�k4�)�9n��'C.����n�h�Ւ=L;{�}�2����yK.y����&Jȏ�����C<v%ĈJݦ��ź
����~�p�g�1qRN<�fvk�S������#w�0�e��'(��	�.�}�x��i++�{�>!��.�GHl�h������_8����`�_��l�v��L�^�v��!���W܅1Oy�&�'aށB)�a�5�m$p՜��3��!l)��i7�z��dX��d�ϩGCz)�5ۄ�����^�fj�m�ON���G%7�CW)�dY�֒T�f�C�a`���
o��:_����פ��.��(�O`�yg#��Q����"��D�]-��}���%3�����+�{��m�9q؊`Z֛���6�m�N�]�vDsr�y˔�����3�`�M�>c<(D�7/c�)j���O�����k���m��:w��������wb�1k�x��$r���h���*���&������O��A��Ɍ�ֹ�q#�q�>�h˸��5���	2�M!�"�6�Z?za��>��z4�|?\��y��~0�'�w��e���'�U�u0��6�5ot0}�?�PBZ8D�4�3đA���7�B&2��3�Z�o�S�
0=�Z0'���||��ѡ��]S�\��"���7�,}v�]�x�j̸�`G�4�H*��`$]s�4$�;�r��g�Xh,�ڊ����ubU"�]�M� �
eCN�����}2���fxK՗-@MߙNsP��>r�]��<>�;~�7nvȊW��ټcN��b�䲱u��r��{�����I%%�/�23	�@�R��P��/��
0�b�����1�?��QP��{Y��������aşs��h�j�2�q;/:&��L"XT���<�8�~�����4T- �t,гx���G4�Z�+}�-���d��(��T�O���Br�3V�(�%�Up�@#e?z���,�o#�ݳw.��x�z�.=[D[�݁��$�A��-�Yr��O��>������8�~y��1��k%"a���������,�����+߳Ng��Hb3���M�M�x��X
i��:�m{�'��QT֌�il)��^��>�m�\نg~|d|�s{�8[�ךQ��x����A���G!�+چ���s�	^�+�.'8�ת��`�n"O�il�Y��(&�m���_jP�&�ߕ��gJSλ>��p\�:&l'�F�6a@ o2�!��A��.����`P�-�r$�z=�/G ć�L���w��8���Y�bX>D�6N�����,�z��|��ms��>��+\��ܟ�������l�_n�7��Kg���|�4h��_����|��iT�m/ HK�:XH��i����bn.v��g�[ՐF�����v�j�җP�δ�ۑg���w+�@z}Е|��m�2�~qQ�%�|��Pqɦ��#g�*</�t n}�k�~�f�rWz�N�Uw�.�
���kH1Û�Q\�g�M����0>OX�z��f����!�ټ���V�7Y�XUQ��JT�I5cE�×��l��#��7���&32Pm�]�¥�ޟ� �"w���*�?_l-�7�̕-������:�L�"`R�mv/�f�\}�@�m?şM���/�����o�t?e@O�M�"{�&�A�S�O��~&���8�2�&0} �c^�Q���ɚ�
7�/��gr��+jQ����~z�%H��U:��hS�":LH�l+�-K�X:DX�M�
8�{���[V��`9D,ە�k�N�|�(��%�UIyo��Y�.��"14U�K��'�}�̖X�IӸ�*-N�冨E�z����0�d�����ǥ����$�GZ���������$�`Rjk���L�����v���\|w��"�3�侙��U��Hm�mص�M�����95"\�:�K<I��QZܲ���+��rDa{�����h�)��掌�Y�!�@���a�Y��-w�������>n�b)>�X�T��S|{ٗbN�ZQ��		y�ۀ�@%���>���z61���J�Vh3V�w��a�%	�͉EDr��Usp�uxQj)�Xr�F��oBA�|�"ut�s&>�_���YVP!��(��#z��KZ4t�����t뤻��'@�Ϗ�/u�x���ZJ&��_��3K��f Tm�o9M*�^E0�Ό�o&�i�^�Y36:)���N���Xfڃ2������}׳��'Q�}�j���#iɃ|�}8	�\&��a �1q��8�����rj�z2�E�|>�K!Efz�,�	V=O����P�7pE3G)�����Y�� Bg
M|�9�:��ɐS8c��q�mI<Y�<=UG�y���4���/7�b��;���Պ����e��i�;�.��+�_��W����5K{T���O3^qwӮi�; �Q/����F`�[��i#���3��M���v��}�[��3�e�tR�K���g�\�w%����h�1�vA����-��qGA&	0=��/�D+w�.�����E�P�[xry4	��(i[^�R~�|Vq��+$L��
��h�3�n�Ŷ9Wc&�l JS�9���D7/5�S�!�فڛ�@Z��;�}��hb���׶�	�V/��ܮ�fnco�yK�;�v05鴽�<<��`T=���	6u��"�ì���Nli����X%gpN���<�}z(�U?�eN�3D����S�	���tQIK�����'���u$ؤ�l�)9��T��i�vKm�M������a`kg?�gR�b��1>Fa�ej��'ٔ�f��:�ɴ�p5��7}^Q��r��hWmN(����!�z��j�x₌X�n�j��t|��RcϬ�r��kML�*L�ِ�%�K��*��LFr�=0i�82$�}� �����g�Q,7�#��o��ۘ�����Ο�h�uC_��ח��*G�'
�X��U�V��@O��}:e�);ڀeC����K��1�E��S�fjuG��OS'T��R}����W��2��'Ŗ,�*n{jѷ��i���(-ia��4>+(��p��O+�Ц�Ad��2��
�&b�,�g�w�Vٝ��@�7k�#?��DmOxb��b�r�H`I�+�'��(�ږ��.�s�9oYS+=�N�oIR���Qĩze*ݼ����$�����|��+�K�ϱ��^h��������/>S���Z~qq<{�)��2I�XC0��E���Bz�����SM\oh�F:x��͍bXՙe!cS29T17ߘ�<�۽C�Y��P�Zc�1��?�d�I�J�9c���]O�+~�]�i��ϰ�>�KD������T|�b�ӏɋV�����c�_�+�~9YmT�a��8{��ͦԤ�t�<��d��9��}9R�,lx�Zyy�P٪�������3,}��-A7!�g��� �'��̩�eA�����P1�V�^���s�,.�iZg�oX�;��c��azmN�y�z6���Ϭ�?>m��A���A�^�mH�q"0���-�5����.�DHm7(���g�v��盕���s8����~0xg	�@e����'�*m�B6/9��!���v�˰0S�t�����G��i6qM>��<_��d�$����s�,�������M�F\[u �C�WD��)'=g�����
S��j��S� ���Hc12�P!ώ/��	�Oz4�ش<��)���ݼno�LV�[��ѐD}��h���&�k�/te���O=�����5�I��-{�Kr�l����{�>�t��8�)����3,Ûz�/\3%�	���X/��16").�֋2fjE���篟���Yؐ^��I�B�/۝����+.��֔�������d �B�����}fd?�b�SN�Ǚ<�C$��|kT�3;plPt�c�K�*;�uKӚ� (��N*˵�}sE�y's�&$^������a	��8��_�+��r�u�=��䁟�[�+`��_/lUk��H����3nfGB��Y��x�s�m�I)���n�i=�Bj<��u�2�Wxc�a6i��~���|� ��3�9����/��1_NWQ�q�6���pho�=���P��O�L����"	��| :�m�'���"K�'Pi(��23�%1�̑�7�U�"Z�/L�oh`"]<Д��i�1�f&CRx��z�%�zo�]r��6��H:�e}�TPl��%׽�L���{�on���fX��G��{�N�f�.�\�qC�,�[09�%���{�7(��Mcz(V�5�E���� 7K������q�J�T�|A��S��3ea�$q)�� rA����D� $M� C��:�6��ͬ0a�&����]�
aRLa���
2C�_Y��}UY�M�.�A������{�����[��*��1/�O\"��v��3�rL�e��^���O3�<[F[��[؝�VT�us��6!��(	@n�MlP��0>S��ݻ������d��F-���Y��ݪ��i��M��]u���f�i�T��|�\�ް����� ����
v���������c�A�
q*KAe��z�v�f�&����/�̍��BJ��~tz�"^8�޷�.X�����Uژ�?�ᨉ���"�$�ބ��
��+r=�_��_>�锏��g�0���X�vG�l��z�+ {�rG;��~�vu'=���eƞi��Ԗ��'Ŏ��,/C�����B��W�-��+ ���z����~��5�6=)jn�J,m��r�u���M=�D"�x�yq��#��x�w�!�zQ]�j��'�G@Ncs��+ $�_��I-�SZ��Q�0M��~?=��Pʝ�(�f�ݙU阘�tb�,���e���P��@���i�]��h��&{Ȯ�<4#/־��W��vsT��He��TU&E��u��$�%~zgH����P?�T��h��aI��!���7��XQ�`���'����X|Y��'�׵@,mH��|��|��oa�ȻO����n��=�̸���j��Ե|\7/�p�7�Dl��=��f��V�"ps/U�3�*�ƴex|xh;q�hI|Y ���9��hP>���4�O#eh8	�yI�x�?R(��������e4��uR��{X�?-D5)^�r�nj��&�V�m崓�z�Ǐ�F=�՘W��H��WTNǮ7r>�	ň�����wئ�&��qY�ѩ�� 8�m4�	>��Bg��\F�)�ʺ^Md1�e1@�`�y.�Vg=������m鞚db�M,��{W2��r�T����)��zhץ�m�+f�,>~S#(��(�xV|�/yL|`�ۛ��I̓��>�&Q���3Ł�:��Z ٣Ɓ-�����Y�1ā�������`�
��vJ���L�VH�c�(��^4��L�eO���0����^G�	�)�(q!,x2+&+M�e\К�R@p\��=��A*/��PEW��|��n�V��	h���$wDy�R&/I+	&��Yj2#�7�c����ղ�p������8;EV��o�4�k�_1\�R �=1��n�9���ۚ���A��&�ae��(��̍�������ḧ�Kx�%��~v�B� ���ǃ+?3�֠�S����	C��a���p����!v�]妣�s���τZ�g�2��$7�2�]{n�/c�qe�qx^���j���Dc�߭!��5{l�r��q~��a��9v��� ƖA~w���C���p���ܧH�sc�����!�M��Q1������%9K�RZ,$���q�q�+�J�K�R!�F�/��m��[3���XiM�ZLX���q��Y�����vlߣ����*_h-m!s�x�"��	�`gR�}�`ZYx��2�'��.c)��F�B֎�����b=�-yA뙛�X�����U����x��%�A+��3 \IcP:D�%�܍�YF����?شS>�$�N�
yQ�,ӅT������-֕ʠ�������G�,ǌa�a6~��k}E�&�	��NJ�ˆ��<���⊃a�xK�\������L��s����QJ�on�g2��u�N�����&���/cU4¼� ާ�횉�Q,%X%�����?��}��	X�dW�����&�l�5l�o�f�TD']�T�(����qǎ$)����D��Ƨ�Z`7��� 3�Q2�jB3���d�e��e�<�G������c����Y��wAcj���O�$qL7�a�ye!Ko	oo������g��CO��`�H���*C�p���D#��"�/,k��x�Վ�P��YOؾj�}ѥC��vC�Y0q1#���f"���0l�D�Q�3�P1���g�ڠE��N�+�wSŃ�KD��� ��v�PxK4�P��s\+��?�ʃ摮�&�C�Ո�F�]Yl���L�l:8���[B7���κ�uߚUR|��q��~d�1�=6�A� +7��8��3�U1���O�Dܡr"�z�jm� (]<�IӋj�!�`߀�����ڽ��é(�������촿@W΅��+`g�ű}A_�iM�;�s���<�V���t���!)�,�X�����a%���[y����l��cΒ��Aa��.��~U�����SUp��4����ߌ�QKCS8k���ef�y-�+r�M#TR~����=��&�(�����p����BQ�
�q���P4����z	|�ó�ξ9�Y�=z�kHJL�X���� ��hq����Q+������9����#yF�����R�z`Ϊ`��at�߁������ы��u��ү��Ag}׿���\	'��*C���DN����H~��߻ѵ��#}��-w\g���g����|����(p�(�H={��Ҹ_�(an�h��[MSG<ҡ�%�7�;k�����'��\.2*� 0T�y�F��4E��
HR�]ڜ8������)���I-���zp��a�R���ьGF��b���(�a�aH�yڝ`L���Լ�X��`���e����&��ӏ�c�/�A�Q�dgyM?*e|M���'��?h�/�m���Ul�����?��M���moN`���Q��9?7�0:*���U��f�O�v�j#s����o~��������[�����z���b6�$��&xJlZɛQ&��a�O1r�5},�����D����G[v�����}lNif�̈vqW��ۀp��v��Gv��쑇�c�7>R���Jk �ܸ�y���M=r�IF�L0+��A߮U�C�{�b,z{������J��"O$�\��irB1�׋t})�g�_.ny�[/�L\䛖��l��iN^� 2,%(�]^�v��P^*�,��e�����-h.t2����%��?�L�Dj�5��-����~s��gݡY{�\�2�`��u�3ύ{灾w�7�:��y�#�����r�>��Q��K�{���9{m�n��fp�Y�D�`��v0ɗp�6ˏ�%�q1O�����`�Ho39�Vh�S�*^�}	a6d��S��N/1����l�#�4�4"H`)my�ר�O�^��gK��pCP� $�[�lQ�m�����\m�p�a;�%V��WRd���or��6�Dӿ����f��>%�VA͋g��E�T��&���e<��޶_�(�����j�~��Vq�*w����뽿��+M�}.~�2l�2z|�
�9�~�OIR{�z>�k�'ؼ�:�vs���W�I���2�$��"�fSχ������ƛ��Q�k�0ޅα�o;�,��R�,�T�C���T*����ec�KI�s:<O1��a��LWV(VEEt=��%�T���܃�3/��be+#�������q��}�s��=�5�Ø�P�p�aj�B�!��kct�B�KVbN׫_��.l�M����H�xh�H"Q0��^�᳃ñ�� o��v�%ڀ�G�n���w�5�܉�u���B?+�a��w�Ⱦ�FϪ׿K8�#70�,��/������n��6��������#Q�d��PW��;�R�%X��?�W�'�qO�ȼS��ܚ#؋GɱY�fO�Pw�}��z�xy�rW��8�Lr�!4�������6a�5�{�Y8���F~�!���S�y�(e/�H���{�T'���Kq���X��h+כm/����zYfs�\��,@�}�"������)�ݸ�����E�@q$���Ț�Xl���n[�l�T*�jұ�?�6�ҫl�,�۟���!��a�V]!������ �5o~�^��$��s�W@%�bO����1GMǛ���Fl���9�Wrb[����B�464WҴю��.ʲ�G��q����}�U�~��] �&��~�F�Lz]ț�6�b�7�J�]^K��c�+h[��F�U}w5x?CЦ�0���G.D�Ye��|k�ĺ�!u�������vzx�S/�ӆ�z���#]��qO�*T^����d�Zʾ$!Hi�����L]��\��@�7uW�����qX�+�fLQ��E��y��C�����J���	=F�R�H��1<S�dxd�H�[�^�7�BTDKS��J�#�����d]e��[�-� ��ؤ��c)G3��'��%G6E�$mJC���KĨ%�=��)jG�n4�؈4��4��%�Qo���pѭ���	��|%�O?�Y)�G_��u�ҽ2�[x���S�K���+@&�tWfI|�����e=Fg���b�~]��{���t��ũ��n�;ŗ'�?\$���?����2��2%��2���]����F�#�_���6T���p��Q���܊#��=n�dU<��{p��������wI_@� �o����2݅�Q,�å4b	�:KE~�G��"�����9c�r��
D�9x'��}j�����W�oK�G �M-�I �R>P�2z�.iN"��_n��吒9\��v�$��"qO�E�bݤ���ô3�N��b})�aR&��
l�ՠ�oL�ض	�#�eJ��1ƻ������爇~���*]
�%���ȝV���cèi����8�6	Md�-�{)��&�{�H�2��c����Hԩ�}Η"����3�Ƿ�q�`_1C��_��� �!�Q���f��Fݵp�H#]).p;�@У�~L�H�Ϻig��\	"i�{	b8��'�_F�]?�>��A���"Qg$�hP�\ς��j�/��	������b��N��s���ppw~���qٻDS7�{0���V�=����𫐷�k��)���F;38n�y-��dS���3<�S"Y� w)*�d�8����\D�y������.���Y�Sm�Tܠ���?p�Ƥ�c D�������\������P�5��N��\�\A]�ީL7^Sjn�W�`0���� 9�S��Џ"�\����!�-'�'�X`�ͫ��0M�WHLp�C#Ad3�D�b�R1�T��D��D���٦H����}U[���y��ɥ�R>�������0(��~l@u]�N#l3��� 1GHΊ=���cZ��S%��_�W���~���'��zm��[~��U��x鵟�IŲ��S3�{�z8��e�œ����%���N���� ϰ�����}��F���X��8���B{V�SØR�tۨ����}�zԽ('$�ʭlJ��p���]�h5�r���K:���i8='���5�G���r��.��#ޢ��˴�}(�"k�2[�t,�4�-��g��7b���w���!�y/��3^XbDS���t8���l��li�Y^��\���K�JG��\�C��+��q��:u�͠��JK�T�*�֨�$;��;��"��K̑+I�o7<ln���E�%T�&&#J���$}���`��pOĝ�·!xl_{`0L���6���h� ���_�6U�{$h�����A�8'���$V���w�64]*�ze��!�)��h��nk`����7b5��8������N,�9=`�x����w����8p�.����M���x����F��ا�ڢF�I7��ʡ�9.�Xso�wi�!�T� ��O����*�}<�T�L��	&d/��FM'�'���"�W	� ��C�y_� ���?�� �ˆFqy,ô�T��i�M3��Y?o����`�}1�Z�~%b0�_"J��.�/fgs��q���/f� JSU��5�q��ԣԲZ��8J��?c���i�
�9J.r�c��Xj(�4x
&Ҫ��[{l�u���X"��ϭ�.�h��W ��z�Dp�=�kZǚ���oc/�Α�e���_p|��(�x̞P�{�HJT���}6�{�,����6�Z�㻝��\���Տ<�s݅Dw��Lx������\K!�5$������ܜ�z�ʾ�%<Ф�]E�T#g�p��k>�
��1�&<׻&�������Y����7��3?G�2�6�����$B�}�;� ��H���O�;�<>��Q\A{�ҴA]?�,Nv}"ZV�w��P��PF�BdH0$��t̍*��ޞn����e4n��E�s����d[�6)�\S��r-�����TF\"���S	t�?3��[����K}
�q?��$�CX���5��6��r<OB$�V`:�B�_�/f6@�-���'�QA[kG-��;ᦋ�j�׺�o�R��%M�t�7����G��� i ���+�(S!����'qIbq?���mg����Q.���V.�J�`��S��ƻ�c�%���!���bO6�*�[��.|#���B'�z�e�i�/G|�K���R_���лB���R�0{�9k���g����&$�#h��X�	����(�i`�@M��//��B�4�Z��@���4�>�ԥ��O�k��M�M����{*�&84���7#'aj���������d�R�(�����r�Pa��^�x��k�ω`�.���~aH�z�W��;>F���YM�'n����B%ˠQ�b��wȕ��"��U���A�%�5�?=:^�g���֐�ʤV��b��=��O���������&���v�/�ũp�=,�Pl-�,�c�$�\
nKJI:�`��K�o_ҳnE-m��]���\�S��Qm�T���>��(`Ro5�q����y&�=6��Z"۬_- �\����_<s��,*#>$�	�?f�/����ȿ9[�[��J��Գ@�o�f����w�d�A��Fm8,��Q�x��� �!���h�&Mȧ������Zl�z�`��tE�����P�ϭ�o�7�w������@UJ
jvW�]*jD�T*����A.+��5�EWWLn���������I��MIPҫ��_����L��Sƛ����@��;f?|�x���~���N�e�~2���ȏg�ʾխRT����� 2��%��z^�5h�#�پ��/
T�z5�?�?��NW�'��4���A6����ǁ��E�Cy1L:
1��E��c�%GM~P��s�5L����ɓP�F�@G�y�&m��vh6!���c��f� %�Km��� W*t1r����rb��칢M~m���P	���m�����!iM �M����p�n
=��ɍo1x���T% �����c�K�i�����3��X�d��;��H���:iP�ŕ.ԫ�������M�G"��e�.�Uw�QP�:�Wf�a�g�`��躸l�r�L ,�W�ܓ�$ !5�CQ.��qU~6�3PV�$����3�O�Wl���-���������iWQeoߞ�K�����(:�)E\%�$R�~� �da������m�xZT��PN&�|�UZX��o�T�xi�G���ʠ����u�Ct�o-+v�O*ͷ�J��I��=m:sd�E�56����D�'�h*!}�J�ϺiM(fY��M�����«M]���q3*$���y{��8k��$�Og!8����x}$���K����}tK��6�L��b6�MK̐\T�����.�X�U���ƣ3<$�2�}w騡Y<^� ގnPW�D\�m3�Q�no�ʡM��
F�̘�qN.ޕE�ࠜ_�Ɲy�Oh@�oK8�y�TĴoi��l{F�\�L#�������G;(�{θ��;�	��!	H�����2�W��m����^�z��O����ZV	(�Na�)l>g�I����B��<���?��=�y؁���[�w�$��Y����
�<QAXI-����`8㳨�fJ���0��������M9⦴�����,�ڇQ4�m|]B���,��:HR�smC�q��U�'��V���1�I(rզ��HǙ�)�*[6��7�܇ᾟ	e��;���𳚲=�3o��B;�DBy65|�MXrumt�%洫���=���M��EL�1D{�Ep�y9T��&�hU-���휉�~��S��]��m�n���d���w�e�q���i.��ZC��F��⤑<�1�r��
Q�N|⢔6�Z�8��gf�鱒�μCvya�Z�"�:l��z��d��wV��I>��8`G�g�1��~��򔥤����o��^�:3� ���Ye�����MjԶ��J�A]�ͯ]x���[=��_ݟb�H�_��	_���"��5�E�w��n6jө��M\�>�(꾞��"&2��D�!+�t�)��-V�T��+ ;%M��l�C,^\�����_'`�,�%��	�J��Ư�[x���W;�iL0D�j�6�Q(^v���5�Ղ8I��Fݦ>8��ADF;�^�a@;9+C��\���RU	����
�~P܆��$���u�!#�aN�`ņ���^�3���M���e'��3_�<y����A�&�_�~�\����S�w�7a�wB�K�/]���{�S]\Wt�:�;�����T��w�]�����36��Z`fc:��`­���.
y���Vt����+;����]+��*/��G3�n�w|J|h�Ķ�թ~9�����q�;�ԍ�NvSZ
��_���Y/��R�;� @��ώB����+d��/E�3�x���d�8�����"��Ct�9f���5"0{~���8��N�w ��/t���xu:ڞW<~�����!Y�8�f��31���5Eg<�H�i,�l<���5jb�*;Xo�ѷ���d"��F�jv��?E
�zta���7��;݃�KC����$e�m:�\�!ө\�=_����q���v��T�<V,ތj��0�&�H�4N�0�ʟ��QA�E%F�ك��r?Ėy�_1;)�&|œ恳`7L73}r�m����6�9���),���Y
(�%� >h�Ԅ��w�|1KZ��c�y_ү�79�Iz'���/8�f  � ������sR�9>�ߺ܅,Y��_o�5,&o%�Cۓ��}4��+B���|iX���f�ه�܀C4s͜$�Pu�� ����Q�z���Ã��_��H��XNVd67�jG�1�6C�s0���9�l��+ ���_��_�,�$�s�l�Y�`%Ð����ر9�b�m���n�l�׻�L���_��Ϧg*~Q*_��l�=�p,��t��&�,�w�.O�����q��vާQ�\I�a�E4<%%:�k����g3*8��̂��S[-v�o6���ogx���;럨�+�
��i�@ctԚ�n<�)[!QJ�`��ٛeg�/�r���ȕڊ�I����b齹�ә?���;���h����̍Y�i�}��|,���N�\� R��4�?��Y�����HI��x��0��[TԶ��٩�(�]�;����	��Ō��b�i�A����"#��[�0����	����t03PT�u���]�ʧ�ߖ[�i��6�5�%���I���"B�u���{�C;����I��:��xi�N�40ߜd����.׭�|���A�5/csd�j�����t�~��H6�=�7I�l*Pw�*ӆ&P�O)QI4���<�����!g~�9�wgK��߳
���������)��Gc>Ӈ�Y/�|P㌡���ܣ]]��Å^�2�**�T��@?�c��Fbk��(?>�iϱ����"��/�ŝXAH/ny�m_�D,x�Zp���{��tO;k�`�28��H�B�*���7�8S��*D]�&�W�힖�c��F��Oq*\��pD��n҇`�u*����saMnq��H���g�tY:
��d#H�l�o����`xsM:~�nD���
NG���G�����UM��Dg�`��G&�b�T�K�	�0k;�)-�)��3�U��i���8>�9}F�\�5��}���yz��i�?
,��q���t�p�f��
���jͮ}kA�� �iN��R9�1�'o�B+S��O�Z�͚D:�?��W��O$N:R�B� �
%��/E���vt��������� �3uJ��3�^Vv���w,&��`�Ja`ƪ�q6��;��iru��ٞ�����z/ �U���M��/��9$59�4�$�ܔbB��rE��t��1���0���d�s�
#�C�����&�&�T1�!IO;���~X1m_�^d�3iF�!��z��O8j��Ƈ6��lu�瓵���e���4�\��"���4x�q_I)���<>��w^���g!2����_N����j�hJ 5��^y�!��¥e$fȉF9�\�� ���w�����4?ǟ�H_ՉԴ�� nMϋ��`�!��$�j��_�He��w5L#��"^zĭ�TA�&Ʒ =,�~����4��m�^�9�ȩ)lv����|0��	�iŷ��HQ�Y��3�O�����8�����2�J�OI�.�.&�Y
�ah���e6�V��x���e!��4��b�L���n�G���?�%�%�T����ϫ��OS@"#�O�f�y�ӵt�ď��H������%�,���#�h����=����_���0�
��|��c! ��o � ��CL��+.��k�l����;XA��w�>��m���Q�;�Z�~�p@�¿�oڵ�e�Q��x�%ǉ�����^�H���ψ�xZX��Mj�ѸݕrC?��C�NvX�qvL��?�"\.�'e�E�呛�CIE���(Y�:i)]���z�M<�e�z�4ߋ4����\��? !@޿����xZ��C���O>� �\�.�Ǿ�������B�^_�����u.��|�.�&�﨡�/��\5��ݹݐ�G��2�۴���]����ѿ̫5g.��M��z������|��&�.�i���s��.ͬ���?<�����-���'�q�䩟�g���j�k��:���NY��a�^m�Gk�l�|9ֶ`��;���ļ����s5f���#P �}Y���V��X�o��5����ߌO2�O�ϗ�����ߺ���������t�͑� �#���@���-��Y��M�\� S�9���� ���/�,C�[׸\���)�>Mϙf|�ō�5)*�ʗr�"L�x��Z>Rc �:�b>_��n���/uTt祛T�)U�툆�9,��Q�iƿ�w<�h���-C�1x)�j�|}�_d�V6�~K�%�]�X��� }o�W� �����5��χNq���)k���׉D��)�Z7��7�M���l��_�+>����Ý��>b$�� ��k|��`/��W�3ogTד������-5�~�;���Z�����nI��I�P�+�_��)���K·z�5��7鷙e�k��ӕ���*���]����}��ٿ�ЅT0�>/�����X�"̹�[���(x�y��LfQ�K�q^�KGei��T���y˿��t��Q����MVW�����j**����_��\�ղ�y�+f�z~?��	ܻ��o>a��kJ�>� ƌx�WQ��>��%��W��W�E>����U�x�
�]�Ŭ�I/�� d�Z�2Ԍ�'���^%ҭ�J�@)n�ny� !K�A�񉉈Ο�Y�
v���D�59�ʲ�mVJP �XI@Tb�W�D���G�#w<�6��SWL�U�s�Je��:��sGv�:/�l:�_�|g�+3}v���;����ȾN�-��2xe[1yf�w6%C妼[��*2)4q����p�����p@A��Ƌy�q�v�S��/P�7�/�ic�c[|D[�S��$�]��*�/6�A�w���c?�;4�X5 m0�Q%�!c��Tn��z#F��A<���������!>b��E$�NfoX�A��*2��z.��/����?�8���v���5�G��Tֻ?�ı�@}�����CIi��V+[�j�N�9E4�9F��a�����Xah����!e��ؖS�/~gŕ�/>[6,����O����z&?�o1h�)��������?B�>7kA*���1 [���|�M�9<�c\Kx
^�Y��(B:�S�^&�#,7�.�lT�I��g���T�XY�
h9�����Ks��n�l��_̵��P�zI�YC7Ia�|A3�wD#��\�}���4�^&qZn�Ɉ�q�4f�8�r��FsN"�����f���K�sF�<D���`��L�ڵ�4�CT�ז��a���3��z��H�ש�3�f�&r����Ed����NZ��=@�	�΄��J�d�����VGV���]y�����[��D��m�+A�����& V
�����Pʡ@ 6��9��
�ƕ���s���	GZ,�wVїMj+��v ��r��C�n��L��������z��R��p)ðƄ�%�2�}`���F��:v`4`8���R���Pex}W0�F1%5����� ��Ԣ�"K�q��wW�w_h��X�)��J��bY�8��%���!s�4����w%U���x�M��R��!̱6�r��D"�Z�>��$b�Ie�}A0˾�H�n�[a���d���l3��L�\
�,Pj�����}El�4f��D����cxo1�/����X1KQ�|**�&"���b�E*�kz�b�uo�1(��#5@.-�~�@��|����\�T��/!&�_z@���P  
��'p'P��ճ���Jea�)E�il���dil�U�6l��{g��k�� �[m#���q+WIxn�t��l���[x}�����}��~M��BA��`�Уt8��\M�[�T��ѢU�Ջ,=s��v�����K�qN&F�*8�t�'@����`W�Za���9v���Il�cܼN*\��{����[R���٨}�a���	mx7�ܣ����N�Ȗ�d4�Ր��0?�y�s H���e�G[�L�8i�)�F���ڮ�[��1�z`�:��X�N
]'ܭ�����V�E����wߚ��P��� isF�W��s�8���5�<��J�1G��s�[�X�	K��K�� �ߋ��,�4Lu1S���c�j��"<��怱Iub�$,B�8��}�=�sk-�<� ^�k�>}Gܨ�#U��_��w�r+<�[�g<��R<�w�B�	�"�i/}��kW��t_��6��/4K٫�a�T���.c���@%-;g1F�� �-!1ã�2�0���z'~nR�@�f	o���`B�f$_Vj�:��#���V�)�Yk�(PUH���Z�d���j��S �Y���hv1ķ�V6_]�r�'�Q����������V�?�.:F&(��jm��2����!)|��ӗʚ̺N��DB�>(#�>m'U��gǸ;��ی�U��J����+�R�����e	�c3��?�*ʗ������^��+ȭ���[k���)�����48��`�k*��;�W!����U�;U�D�y�a�1�_�5�֪{��(�B�!�AOd�|Z����.<�c>`�5�����]^�]r���+�����!�+�-j	©��!��Qg*R�<x�,�(Y
�w����u�!�A��	��iK��%6�-�������ҵ�r�K�����v�Lz�%�ӥ�)�Z�ң ]ڏT ep"s�E�u�d�eM���w\B4�����%�` ��_(�+�V���v�VW;�k�d�K�_G�Mj�U���[1P@^St6��*�Nۏ+JvpD�J�ڽ#0o]���0�:%�t)����gdo�	�j���P^�P`�d��G�'����gՒ�-�E��Ň�1ջ�X�{k�$���)h/r*�h��(�U(+_��^��F]��q�T��V���� ��T8Չ���_1{��\'��x�+ee��D������`���;� �3��N�����F�"�]�99���"ܘJ#>k#ȷ��U��v�eu����E�� /�s�V� ��iP�n3pt�
]��|�����<�Y��g���hp��Q�>`5X�f`A���K�a\TԜ3P�h�÷��4vesjmM�UK�J�7o� Q}%�^���pu.��/r\��1��ړ��#�t�GPY�^Lю��w��e�?�G\��<��� ��A�����b�dQc6���8W�w"�#��b+ȑ� 쾨�F�Вx	_M\ \јU �ʪ�qB~y��w����{te>f���R�]��U2Q�����r��� .���s�֠a��V�':�
[�m1�z�/��x^|p�*�����r��a��;�[�7��?������(gE������QϹ��d�%� _.%4l�{�,yט-�'��y�D�{���Gk�J��q
ʀ��.��~#ay�Ej������R�GѠ�f�<���z�n�3/�0LT��m�n�1��Li�	R����8-�0Lm�Zx%���B,'4B:խ8��P{oL��$�8?ӄbJ;Z)�OX{:b��4A�\�T���ٹP�R��[`I|������A�%%?a��U�w�L�Zi�Fw��l��9��(����*n GEsy=�S)�]F;n��ͼ\h����J������2s{��뤳��µ��ܱ�i�7����l��c��!:���}Љɞ���<TG�Y2��Es2�@z\da}� (�����S3��=��/ԫ<]�BE���`h�G��6F��Vɫ���*d��W���V]��a�`����cP����E�6�;�y���\�4<�˪4�W���a���&4Z!�)�2
�<��	
e��^.�B�P�1���u��]��x����G|�MqϽ�j�	C��@�"�:|JQ9�-�}��N
��s� 2��/��������:s��� 	pA��"������J��5ܬ�}�Wj���A�~O;��<�W�縟Ͽ���[��[�~f.4L�V~`���0~gv�Kb	X~�%k*�Q]_Q����Ja���{�j`3���)����]���DA�\�� +�@�Z��~|�ݮ9����GT�?�xcx�����B��S_���͐O����Y矶<��	�����"�)���j!Mխ��ӯS(!Ī�o���8�f</�0T0^;�B(���3��P�;����
n��Ѣ7��x�Qgy���N;����F������H�+���Z���w���b?s ���O,�~c���^۩�p���[I�lͼJۊjK��p�g0{�L�M��fm���V�f`Ә&�s3�L���ʡ����+n��/����~#o��2�x�j-�G�Y��aI�Zե���(�6����b{e˃��9���}��F��/���>�3�|�}�c9�x��mw�{`�5�Eݡ<��"�fs�M��G�KlVcs(0���2�ޣo1᝵*�6Ʀځ��Lnw�5���1� 5�>Q� 5���7ޥ�����X⭲�h�6	z ��4�I���<�LK8?��+��o�ɪԋ.��Դ�U��3>n?��a��@]�k�����*�������=�v{�'M�e�w ��GJs�D�6_-�>&ګ���|�,� 0��Cw~q*d~�2۸�2M�ҽ!>g�G3�tgpM�ψ����U�9��S�w��
�y��-��E�2g(���g3�q�:��.���)gq�U�R���33��]E ������U�x����Zs�%,����q�v��c��.��Mtg���SC�3�l�=\d���)1w�˔�ܰͬ�|���\�����\E��q�L��ڲ�i��1��v���/)Db��ø�j�nXҭ���S���$e�V/���\�\��o�L���k�e����d;�d��P�{�� ���o��py�Z�+T4_���ګs�g�?��7)Bܝ�<NL�m�s�%M��|Ά=�˙�,toZ=�C�ל��.��������S���]�� T�[{�/�rߜ����%��������d�[�B���l�ɸ�r�1c��=�;�r���f*�f]q�\|�yK�y3�m�ܥ�ĭ�%� �y!q-g٩��̱��+/!,�]6i��D��E%�*�t˜%Sv�� eK@Z.a?��	`��|�y9�:�-����_8v{�����?����-��X>�'��O����� � v�a�q��z����rm�@<���;]�m|�{��75սFB��s�tK��]Z��pAGC���+`n�KSNe���s�-��"\i���Y����|�mEz�'�.����h+P9֞��N�v��by���K��p� �rwR��/��h�夾AFc���g�����	��s~Χ�����&Z�,Mʐ>底){�Jj_�RƉ�l�k0���Jf�����G�A)}o�:n%���H���`�AU��L�8�q�ޚ�������A�B��2=X79���'��h�I�y*ؼ�	�E� 5��˜�S%o�(���Q�G���,\0�4��:����� p����U�8w���{�l3�=�p�J�3�ODo/�1X�_�Vb^&^v�����0�W�(��������ؤ:�d�`
N*jxW���D������Sj�9�rڒ�p��� �,�Q
S&�{��-���>��R�.V�'9�G���0u���5��x�����9�����b��f�6%� r.5�181�%�Թz����8��`���>��i�ʖ���ֽA����ŧ^r�K)n�%*��~ �WR�߁�m�5�.[\�-f��4��
5R��R.��C�|��pA���Kh���S+y}K���?��x����`�\��#<hoq���'���Qg�����cV�=e��Y��:�^n�����*e䖘�c�x\�®�ȣ%'��@� �9�o��%�`��X��<���5�T"���Fo<���3��]J�R+�v43+�H���F� CBp�r���g�&tr��fS��W�Rm.q3�*b[��Wx�����QG�5��#vbb�x,�@I�n��'> �+k��UZq��Ҝx��:b0�;SBN������a��k %ئ?�<{ ��E��g��6��F���z�By���4=�W���سZ�-��>5����T�+�>����1E��
��*�i�8�1�7EFZ������.Y���s�������������j�r*�M�x��B�_�J�)k���Y̦o�JZ]?��l�������q���&.���������g��Q���.�	��x�91[E� V<�܁���L����Ym�T�5,/,ȷ�\�^����KW����^nx�|����<��T�:�*YcF�1�K�~� O)K��p@��r��G;1N�w|�/>vÂd4�����d���'��YՁ�^�L��/c :������usM�U^c0���_3�Tr�#H��£����� N8����O���j%�r����%�8>鍊���*=:.��|.:M�a�O��b<)u�%<�G���P��T|K�j�b�}j[�������9��^����D���� �SE�p��R+����i�m��/�ϔ��y��'1��jj0\����%�n+0Xl[�*,ձ��M��+눵	m��WZ��%�q�w�r���UŖ�Sk\�*��238s��� f�������2� s�΢̇���Uo�>8�5/���F�u���.j�fz�4���P�f!V2�LK�mQry|�9�ۙl�Y���UbpBw(�?hv|�WW�X`���.%馊w� %��\x�6��Ғ]�|��jg6O��͹���ZK'Ig�`M����.ʊ���N��f|J9�\E� �5��������@UJ�]�f���m���}�--���4��Z�M�B�x*x���S�|�ٗ�� �Pb*C6m�_�5��ؽqǦ���u9�[�Ѳ�7fT�a��_�7�
|�{�M�Kl��,�$uS�%�<�}G� ������~��gP��.�A���`�X\ʛ[�^M�������ؕ���Z�j7� ����a���V�P�G�� ���@}j���w��s���cdy� e��L�X.|�E= Y��q�W�%�뷵^�⿓��y?��IG�*���72�*|��*�S)]fm�%�?��gk$���"O*V&|��� ��-jA��De0�%/�� |�RoN� �U�QϨz�V�(7��7K��d�Qbb��%y�FQ����R}	w7� MˀK������"�t����_�Ds�8{�'9�������T�?勹�=m���1V��q`�4X`���<���P�Vu+P�o��V��a^yȒ�P����y��hm��Q-��0*�m(���rs�������4��UG*���� �e-1i�{u��ͳ�䌳|�>�W�)�y���Td��~& ��w��Zx��}Gf�o"��P�)��Kyb�� �VW�P��"�)W� ;} ����?BV� D��lO��a�)��P��.����/k��T��z���X����o�6��M�mn3t�=�3'�!����� �%kT�E���O��$^E�Ƈ �(�]E%6j��16Ѡ^i��ӆf\�4����Mȗ��K��V^V.z�ڵp�\�J���p2��͘�"3����U瞥��&��A�������O��8�<	�~��A��Q��s[��1n�K�Ħ8ܬ���w� �}����iy��q)��IM���'0 �ŵ�����i������ǫ-���� 0�k�H]�\Z���r\���S�-�Wd�s1�c+��J��J���/
J��y��' T^��l+NB���D\t�����˳�TNӈ�Okg��f�R�-:J׀̙���ɚ����5<��	��@��)U�Y�����a�W��u�W&.�Jw�%��uD�.��ӌ�r����ѳ���ð��:�G�Z�>p����u8%�!L��#�U�e�bZ����KVp�O��w.�p�U�2����Ht���K*Vj Գ��A�2־�T���}l���T��;���'?}L��R�yw=Nv'������Y�`��v'-=����G8��-%��p�e�n�-눍
%s�Yj��o�� +��<E��u���p�W�F8�	�i�p���C�-��_���D��W�T�5�o���>b�a�j�]Qk�ɸ6��cߎ�����x�(�]���&�L�>q(e(B���H� Un���ЍÜ�S�� �/!n�&ҿ����㎢x9\���p��ҎW�c�S"��HZ��ݍuSct��c���]��4ߘ�''��H�P����awx}$����	z�,�K[�u�2y|y�6�\w)EU�s8��|�X㢏�EF�؊)�YI|��?<q*i�g���L����B��D�~���0B�WX��?3cXǙDa�%M���&CA��#7A.l�甙ff�#���0�����Z���3�r�P��9�)�;��f��֏v�>�b�+�����.�H����k�`�x�[h ��u���$�� �k�J{nJ����2�5��_a��XE��qj)bA ,�7�w4:O)J�+%�_;��%yD>�@/x2��ϙ]#��)�nb-9�#�#Prg����8u��
�(�em��0�e�b0.�x^ab�%Ǝ ���x��L5��.L5�d����[�V�Ak$�U�d+4+d�nW�8��m�t߈uB��'��0�/.m`�!倶h�:���A^l���[��H,��Z��8���fUvT ���c��������.�f�G��g��d�7͆?�i��T]�-��6����^L�rJE"�(�8��2�ݵ�'%������[5}�È Va��I�� B�;t5U���a_'Y�o�|ϘN7���`.�V��9��v�S��@`|A�+��7�l�IQ�Ӕ�X߉@�N�)II� � ����W��Y�/қ�"�sAk��'sÉk��S��������%(#B7jG�����LH������Lq�ݗq��5n ��G��+q$�`��
�ළ��D%(9�����ˬm��wT��`g��:�2l�njݧ<ܠإ}x��M�+�SZ�:�:�@8�KrS9�Hx�
?�L�3t����i�L\r7��N".����8��������"�7�F��`�yD���ZW����_��QLx`�����o�"�L0���yu0 �i�0<��q��,3�}�"�n3�XpL�$M���7�n�#�)��Z��_C`��b���?��*X�a��z�x��\�շ�11�|nrx��Fλ�o8eS�{�{�&�,��9�b��joD�bw3]ʹ�DE��0�'_��#B�|����U�d��8i2F���!�^2נv�����pF�v$����{�%-b�ae�f�L�܌! [W9�&��'����qs}ɣb�Ьʑ:� /������Q�0j�au�5��� 50��̝��.ɜ'�]��hx����(|wbõn���J�W<�y؝���ܵ��#fRǩl����7/�)r�譌���ц� S��T��!,2Gc��po�~<��E�<;�m�C潾���&�p��ot�eyY}ƀZ\�)%���6.~�8�㉀��y�n*��/�E��]G'���{����`�F[����B�,�c^ϠF�Ce���k԰6�[og�#ڠ/���Mʞ@���y����Z�}A+��­�1��Zt;����i��X[0�#K�`���D8��*�V>�xRQF3,]���(�QƇA��i��W�����e�쿁5� �\���,��N���A�޾��[��pM��GA�&&��ɟ=�	��̰�7���K����Q�K���<�|_��&�(�jf-�ѯs~sp�r��g�	�6K7)�S �����p:�!] ��U3��;�w.�����������D�5��^��z�R9��c�Xq��*��+��]X:ՙ�Y8e������ ����$Bl�*�
0�R`�C"�=�B|`�Τ��2@�	�ք)j�	����J�W6`]e�.��#�(�9j[�����"��:�S	g��|�lw�b�=�t�c}?V�ˇ���ɿ���p�+}��x�b8�]ͯ�foڅ�g��O�D+R<��c��}� �̌�o��fvm�Z�6��,^nv�E�>�}�I9���h��$�ph�AAf��8P�L2Q9�A2�Ei@%���3ĉ)�n�6���ZH
�M�n�n O�·�;6Ud��9��rpF�
��Rt��mAV]j#ް�*���`ӿ���&��{;�@8���坄���W��
��r6U[��W��� ���1+�}.3�����_T�X�o�V��Z+Ց|y՜ _N)�3�1�n?����R��7�!��5�N�y��[W�^�!�ܹ�%f��,�/i���\F֋��e/KwrW�3S̹i}��,҆�Y��1��/��"R� ��]�"�T9��r��L=�s*�f;�B�ۍH����î�	H9��>YȦ&�(s-��R����Bڬ֡��4)/�Q�F�k�o�\�{���*���k��|��s^����X��bZ��H�K�{���*W��`�C���|�4��i���R[������L�� նc()�����؟S��s�}J	 V��*S�J���F"�*[�z�5��6�x;xeӘh=k���=qW�uΠӕ���:s8�K��k$X��Y�Yu���"]���8��_�?y�Y[4��t8��̏n��K�3�� ���U�Xz˰�q��XNZ�ɿ�Y�,����G𝲵B�<�Fދ6���q���}�lv��B�N��Z��es����|����Q� �����@�i�
�ifvX�M¦t�-���Ϲ.#I�l��䖉[�cK���y2T�W����5�C��a�����nʂK`%��y.����3����Q[����?�/5��ۡ�-����-ӈ��J%X-/���ʯ�p��fe�_��q�AJӃ�t�M�^�@H�@bEچ�E�-�uo&�s�����*`�i
��J�(��m��E�d�VBإ�r�f-�he��a�"9n��2*_�A��~Ȥ�i�5�����Y��ۏ8~�{��&g�p�n ���1�X���:� ���W��}��,f�DKt3c;��q(/����O�U��d-g+��6����N4��;������*	!�ɸ�� ��<�`�;*�%	����� �[���oYhg-�z�Gj��M�W^:f�R�̿�5����<j�>4�8LZP
��x�H�g�o]_�e�NEF��)��.��b/"8H7��v��ҸTe�PJ2��`�P��wL�4��p��}W�1�n_iԶ����Uu��i�9�"Ê��5��B�� �ģ-W�����2��������fL�~�1S�7�A��i�8��0/��^��w��Q���o��� +��)L0������ї����%ܱc`%5sf8��9]ơ������|��$���ľb�NŭA�U�s��nx�w�'� �_oK�� ��k����-X���9�� �x�QP^\��z�8;�-�Ļ�(��lvyf�v�Wiq~�h;Ӹ:;�Ǫ�%����"r�������+^<>������L�~� �jX�iyy8̜��]|��37�\g*e���c7���Bq����̞͙���@��+l����t$~S?�F�~�F�����7��Y��u��3$?�Y��S�`��\��R�Y�Զq�B����#�y/��W�CM���5M�E��Z�s��f�k�t�.� �M�o��ƌ2�h��`����B�d���<ܦ�=��)�q5/ 8J{b�1s�� e0jL��˾R��u���
q}�܃�(c�׉E=��&L���^.ɶ~H��y���s�n��U��]5�~��U�;��.�|���]�f���	mw�Py���|"Usp�8��*�}�"�S�`Ȯ���O2�ݟA�Y���0R�r�C�θ�)���rD�y*j�O����/��iR�w>!?1�~c���_���0�g<��y,���면�(l_��4Z¼J�cžC/�c�rk�_����R�zk��(�A����K�2/�����#��ki��E�'�_=� �F����\���aw,Cl���[�q�
���+{~:���~���J�帽�qi�(��'�'FXs�s)���@9�s� �0�b|��t�FM�?JłS����3.~��{&��"��B?-�0f7)�qxK��Ku36s5W�����4��ܿ�89��{�c������x��Li������>����p.Pq��S�5����k���&y�Te%5K%G�ZHF���2�n��qj\1�_����1��~%��,2��K�s���b���Dmf̗����e��S���pv{  ^�guv�9܌�� Q�~����ܿ�W1��|�@h�(^�=�P��=<_q��lR��PtG��̫a�|߄��ڒ��L��{/�@Kռ�/�ʳ��F��f+]�cN8q*�ǿ:��O?�m��nW�{�U��{�-����:�}nަt��>�o3�}9͚��� S_�Z-be���o��>��kU��Ұ�s,0|~?��/R���_R"��:�0���|�U�B�����}�Ǹo��_$~��Bǡ��vSn�W�;e�L��S�X���=Eݍ!� �[#�=J��Y�� �� �=j����{��xģ����N,���� �N�zbdjG ����c000~3�p��*�Z��������V����sf]�_y�����*ѐV�VNce�LC*���HZ�����3�EHU�f�o�k�R����~q���e�f�(��#2�&�:�툃�,`��� �n�ސ�:"�PE%Ae��TQ(w��U�M�<���l�ߊ�=>�{5�^��� @n��2�mZ����(�h�� �p�ږ�~�0�	(;��a����F�}�p(bd���O6uPF5�<�|���g����V��$�A��eY�'�"�;�P������a�n����'1��{x��5:��2Q����~�F���T��D̬�T&ۻǈ��Uo��K;�hW�޲�8�P���b�\žJ>q;(iN�0�J�Һ��z�������l6c�*���W���q#��S��*=%�!��Z�_O����ڵ+�KmB���A�M�U]ۻ��ʇUWCT�Ģ
��Y���3Bs6���Ĭ*P��G,�Yz�,��!��}8� P1�3����L�;� XD���(B����[0�}���Jϝ�� o@�g[�&y�e�l�
hRY�Li�Yr��h}�r�.���2+�w�K�D�c�u��uA��3M@(�/\8�b) �[����$y����7��r����~����)q��/j���(%�޾!��BW߇=DK���SK���K�nLD6x��ѮI��i|jx�*�iR��&i񿴪r7:�jpj��p/j��ǘa4V��� �^�h�vi��6��g�2�:�A�/��Z�"�X����}ɻ��x)G��}M	��d����n�0��8q�q�}ȵP����I8�4����G�߳�R����+�#xY���29�s�W�/^ �k���G�$l05t�G��t_y�2ݰ�p:���h5�y��]e�K���K$�<AJ���޳͞�pj����.X,Yj��H��O�L)�Oτ����Eu83��^"?H�0��+��}ͯ̠J� 3@c�/���Y�����l�(�9�c��������zKm�q?�@����M��� b`�����u�u�����@�.卡V^�Z$�F���,�9���#$u�[e�R��E��7[ƻ�S֞���S�z1����f�s�2 i�k%Q([.�	+��P�3�,[�1��b���≁~�������� �n������5]\�Z��Q�E���/�C����,�-�P'�E�ޥ�b�P���*X^�vN�i~}B�8�yc�5p�%�̧�2g/u����ďD�p��#e�D���2Z6��Yy����.��C�H�����2���	c��ĽJ��>��R�e�칫�(�E�%�K�O3q���c��{S�d���5f��
�ك�iWF��ܿp�P����ׇ��#�������HϢE��k�-aō��!�Ô�e8�?�J�:�S�����u�2�>"������B��s�7���J�� �량a�xW0.�{��T,�.�� :�O����]B�#�"ז,x�E����
�2��L[���`xy�x����!r���)x�����{�o�d	���ܾ��4M�n��TU�^u����I����C�g���lɡ䉡�Y�N�W��緅J��4�2�&����N�_�"�OAU�ߙ�ԣ��#*QjV���1��ri�Ϯe)��Z�+W�L̩��ԭ[���zķ���5��H��W��k��~���Kn��`&-�K[�)�Ts�,7���2�z�N���u��g��� 1���f��L�.[���U����M�vg�8m�k�3�0���+�7�A����)����t�ԫSao��3^X��O�E������ q��VD��q��<���;&@�L�п�*���� � ���J-�s'�[}��'�>�ih���cY�����wf��5�U�V$���%[�|K�j�{��CI@$� 1*�HE����58�Q$���Vw�}F%����3��=?C1��y��C1�mǉ`��лw��-���*����>�e��
Ռ�t�/��!��k-�`�� %$�"�D$���LR^��5rw)~b�s�|���q��c�a�o�;�)z����p��]���,�4v@��h�-��]-B�S��>eac�Y�{�}�P�q��/� ���W��&g���� �Y�ƾ^���w��JǑt���g�(�S���v�FA�τ���d��Q�����es%$xKǄAy�q(%� ��A��@��΅t�P�E��:�����WB��R�6����9�F������*讯U&��9�B|L�����5y@�\7�1e� b�Y��D�Ƣ�n� Ĥ�/V�����C��'�-YKkn����.n�*a��r6��@f<�Fc����oc,�Ix�x��G�����UB�tǞ(/k9�Q5��K|�!W�Z7�-H�F����(��_to.G�q����N��]}��P��^�֧�C;w��f%Ε<^�U��u��'�?�>8�a�P@\�~z�bb��F�`���,<����lq���0h8q-SG��\u?gdZ��nP�I��nW����~�X!E��PP/9��L�d(+�q��_�1�'pJ��gu�F�}ur���\���xp����4��B9 [vd{�虘�)*y&a��i7��leXCj����>��
d� �b`�W�����X�@�Pu��M[a�r�`U%��px��>��mѡ��[��T��>�@��/{��	�40  �4��JR�e?%�Ơ7Y���&F|!������b%������c�#uRʾl���|ё`�i��O�9;�x���h���7��{��}�F�Qk�����xA'��D���<af�5D9��7s�q/�EW�j����T�e�Mz��Z��*x^h���#�ky]��'"���Th���2*X�i��)ǘ����ts� ٭t.J���q�R�ȼ���z�(��J���Bv�!:��-���|���#��} ]V���7�}��s0�����V=fa��=M�5�3,�ſ��������.SJ/�(�*��Dk��c��B�a��� S�g�">H���KsDϿfl'K���Ù@z_��EݹyJ��_��%��f�ЩBk?�Ĩ�����4��`�I7��)ڷ�F��My�Y%�9�K���q�4b�e�����¸-�:��"Tc�͜�,�����XV�Rs���J�_�y��~�]�Z�XKܸ��J�)��F�~���5�|Kf-�H1�u>�s @�>���Jmܾ��	(kS>�e���ᾃ��i�K#H_6E�U�a35�@wǾ'ɅP����6��8��@S�O��H7���Q;VFNh���4���x�-�������K5wǿZ�_�z��s@4�o^`í�#0Q*�@.;&�U��2��G��%�0km�M A@��o4���z��0d
��)G��T��C�R�ۆ[s<�( ��p��h_� +���1
HN����J��5�r����_�?x73�?�����f��f��@���<97�2�(p������U��|�b�d;��\��ȫ>%))�A.
���k��K������1�h�Ҳ��I�1C��Y���0�	��O�E8:':(WuS�����<q7�֭UG�>���nu��s}�"��׭�a�H����`N*��
;��x"�eY�Pc�U!�eLg}�Es�ܺ�u��h7|�?/���Q�xp��9��*.:��g��;Ty<rtE-���f?�H���#���Q�Ʃ�����j��#Hv\Q�U���ʇNR�r`��0�K[�T�;&iEfч��l[K1�9�^���NL�x�Vg��l����yuy���y_�@�7M�m{JG?��P5�L��+.�����eȮ�A�WKY�w��b��j��̦�#��'�d2ۣ��2�Y�T�( x�j��������;�<�+�?oqiWR̍6�u�q��d���O7a^8�hU��Y�X_���^#:v���=h��u�?��:
t�{���X���V�������"L̈́�F��X��W0z!�e�,�D���'������R��LG��9�!��Lg�e��U��U�V��5��P�?�-b�t9��<��+!�	�|�qW,��_��*֧�_r|S7`&� 0�Y��eI� ��|�+��p��)G	,*Wx�	LT�k��p�G773>�jQ�)5��-l�y�J�)��	�f�r�S���I;�l�pY���ҽ��מ#�^n<�)y1^o�䜏���@��*6l�(v�>�&��CT��V�?3lu�*?�� ^2��&>3�(*��5s`ÔPaɞ	�iJYm���������bc�v��;9%��G��]B���A�����8�-�̼�3��^u7�1�x�(]���e��=�d�����ϗ��~a)�����3�� ś�}UN�#9�`�0�}gY��B�[ebQnĔ���G��f"�E�R��_�r����Wo�^�h����aF���L#��K�������Z�{�J�ZfS��ja�AϏ�����CC)��'F��N�� 'Y��J�AM��p}��`=��p@��P�-����3�Š�s�� �'�Bb*Q��dI��qI��@cf�Ϩ~�r�*�����p���j�*�Y��_Se_A����c��Q^]�)C*��.�C0 T��Fǋ�*p?cI}�L����@PD�� �N�{]�YH�BY��?��`����opwѻ���,��sª6�WP���'��^��.Iu,�7�֢\���0Ky#'8���3���meS�km����5Bߗ��n��;��kY� 7� ɮR��Z���1f�(¹1џR����C�n2=%[w�����r������!+���-��r^��b@2`�s��(���s�
�-��(��<��YI]�
\	��[�-��7ԧ�,�z9a��#:z��C;�E٫��1�ؠ�E���+;հ`���ɸg@��zX�����`��1����O���|Ũ��`��0��'{�J����v��,U��cn��\W��.%�R��@%c�?3R`	�=�|������M�
�/:��P~���Q�T4sm��C%��a�U[�-��+|Ub2�h.�;��Vk�_i����J��m�1*p1Z�����9�������2c��qH������W�P9�2�s{����wy�Ø��Ϙx�D :+J������H����)_�����1#.��w9����4��̩og^:����)V���pI���+���dJ�t�7�6\�u�*���mu�=��(`��ĈM8��}LeҬ���B>���������6���AG��W�2���fe���2����%�q4&)(é���1�w�O�D�n�g@���%�L[|A�S�V#�E�u�g��M�q(jPח�:�/�����y8���}*���o��n��3*58+o?��-�3���Q�����)�q8����)� bXn�j�-7�w��:u����I<.��n�s�Z>�/�9�Bh]l���}�d�5\��P�t��ՖZ�͛�6U�w�y0⛫��l ~t���
u�Lj�a��֎38 Z���7�f�������E{~�%'�����gz?q�vEW��>�� ��{͗�� �B�e/r�Y��,z�*b�Q]�4���V�#��2�����z��%�c���q���ڬ9�rC�|Ď&n������׺�WF�l��M� r!��L��+M��r�pb!G_0eS�]*|K�7v�� ��%B��e����c�#�_r0|Q�AJG�Y���������fR[h=�� �F���}W=�&"O_�3�%$�i�'�)p�Q��Қ���r�3�w'l��˦^QׂYae!���p8`�_�>�&+�W����-�[9�u� ��8B��<u�0å�}�|��4�R���7�=AP�ށ���w%}��ʲ0-}D\F^T{�F�Ʃ<�=1ȟ%���%x��ծ������OA��ߏ��8ɮ��nmh�Y���Ks�c381���ˠ��i.EW�4)4���,�i���I~ �%�q��� G��TVϵ��ۊ� $6׹XB
�W�$y?��8��>\F���]Q ذ�#��[_�v�v�b��U���7��&e��+>���im��L�1�R5�)�_��ʯa]�b��
�0(4͋!w��ф%�o�V!�M)�V�R(m�/��o��0�w���e��u _���_�� DA4����K#��J����
� ��Yw�����_��1ۉ�� ��j�bW�����R��<z�	�ϴ���O�o2�-��3���s̽�ɳ(� B�e�' �O-O�Z�����&���q�ՠ��8��A{�W�)b)�ܤ�#�X��*ߝ�zQ2�,<��,��8m�ů;��83O�q.�=N�y@q|U~�y(�̭�ww�Td�8[����y���B)�Bn(���2^����;�0�gKI��h̵.w��[ �s|���˦Q8�`���]޺���[��[-ky1akz^=^��6�g��zj^�9�Q��Ri���P�0�&KzN��yi�!��J��̩��1�����{�?��%���;8�#N�)_h��Q��»W�9�%�L�1��CaO��o7d9נ���?s΅�_�6��g�1n���:ɗg�l�pwsA:��-��,*��q�m��ʨ�'���v�+w�/B�
ǈ[���ܸR �^�יg^��!�5b�!�v
�m	�7Y�H�S�'���[���������hC��$f�<�J������W�JK�c�Ivr[01�T�ϓ�٘��ߗp�"��r���q��+k������m�y��c��o/��ӓ�&� � �R�n��������&�Z�A����z�� �V!�j�E�c��g��/������Wkz��/P[�CȾӉu�U�U���ex�8c��� npa�6��J���Ծ�ȿR�xq��B���GAO�w��s�U��L!��s}�E�ͅ�:��� `��E�ܺ�dZ�[����:zK��㻅´�?�0L瑀aG#�MT;��6V��2�5�$�ބ�~W;��
��R<Z7�����4�{�3�����p �c�1{~��X%�Ǜ�O����S]�g�(J���s��W��[=~�0���
�O��'�k��7
��H[5_3X����^���`_��6{��::�3�/x|�����z�]��:��C%���_�(����g� �b��C�~�{rB��O��l���0`�F%;��W���f�h���fm~,�^^g.��9���#}��֙�����#�����7�33�K�(cr�S�7�J%p%7�[�h�'�tHC5<W)R��Jy�}[�B�ĥ�&[��^#� �R`���ĭLY�+���wW�.q���X��#������\�1���tC���ܧD9z"/PfīA�z�x�� �3����CGP�ччччч�XGP���>����������>�����      �J`��$H��E ��&�L�� S,^������	�+�_!u1��6�)E�7j�HK�|� �-s��}����h�ft��ڥ��LyA��P�/����۶���`�H$ЫD
|��U�(J�3T�˳ � ���t�^�?EI"��5:�	b��M=��]��v_�Z��B�+��y` ��~��JT(c�R�Ţ k��i�g+���2��B;3��\�e���_�A(�`;M����g��~7��#R�(ȕ�-���L���<a�Cf�e3�할�
l�tR2��ɰ~N�R�!4IJl��D��D� �y� 
l��	�	��e�G�$$���~�p� �M�E�!���0H�z0�@Pl$�e�Y'�:P �V%�t�ym6�%2K���p��#>��C!O�M"�@ ٨�V�ti���;�e�<?�n�M���t�q�$�h��a�f�>_U�@�g��r��� �AJK����7K`������@; )e��1$�T{D��S�AL�b�0� A=�-"�@�IIX-��%��Čy�b��ޯZ}�-0I �L��I�&0��;L!�m K%6I ��"����Tv&�͝!$K� �	�0�0%-ڥ �*�%��}� �I6�E�$p{�n���2.���(� $��Y$6qy��n��u kL�A,0����?f��đ�@� �R!��d�"")4"2�V\��6@�%,�U ��0`2�D*$�����|��0`^1&�  � "ɋ��~I �X�����&�AI��3�9�I &�@h����+�cSNJjxKu��?-B�=g��@j��:�7I��C��Z�K$ 5k A�
��,��&7��|�� d����$�Eh���0Me|���H��F,�Z�^�#_܂L��H�E���@e�xX@�|d�4^h�Hh �	�� �*�~Ԉ�%���`�Z ��	Rx� �x8�g���D�D2Ym�E�HH2��\m�7�}��j=/�H���{("�@b|�p\���3zKy��.
%��խ�pf��F��m6����9�o;���ʁ tH�m<:�߹b�IE��՛��H")x�/;ǽ(a6�����J`ĭ�{�>2�㼲O�t�Y�����8����H�'��|�R��O
uk�P_߰|33�t�l��.	����+�@��Y^��O��<[�l'����zMzA{x|	Ws$"[ "Ӝ�ejnUߜ�-�n�m?���>Q�� �� eV�R�+�b���[|��y'�V\�4��=����1+�|G  �G�$�EQ��&���J�hx�z��#$[	�5�g�肔��ֳ� ���Z����� 4i$D���1V��`F�gj�ȨO+j��o� X��w� :�ŀ.�̺m?$~dM%�mx.^�y�-H�T������or��`��$k	 
v�x�z�tT���$�I �I Q A��+�m�����v�H  �A  ��2�Qb$��#�I  �A$� I��A�$��I @ A �  �I 	     �  @ �  �� +    !1 AQaq������� ��0@P`�� ?�
u%Yx���VPe��>�>v�D�k��������6�ϝ���_�� �3_�]����o�Q)!Ic���CB7�Gh�,i���0�9�q���Yři�7�0�BôX�z�P
�:���h쮯RM��W2 2)����:�Y-3dY"Jl�M84���/��q��Q!�0���3��`��b�!�ϛ��B�#5�x�C�j[� uFb�'8�G��+.ɴ�O#!�u�*	T�B\�ԍP�`W��}���9��\W\�VN8���N����j{��ی�J�V���΂� ��\�iF��_I�7�H��к�o���U˷��I.-����e�7�ԡ�?�iJv�4d��J�-1F�\*�>ɠ�d�s ��p"!p!�����f��oo����*6����6��a�s8�	�od�2j1;�ǝB�
ba��@�Z�T�i��(��q�$��$�1�OiФTZ�o�1;a҄�7a �F�������4�g�D�� �����k�6�H7��v�EBq���CT���Bm�e|{� �� ��s�PR۰���`��t0wO����#?��j�?@%q��h)�L�~��y�%���?�1Q%���ֶ�x���%!t"7��}0��E��0��HrE���6V��)3 H�gl����$l���%d�0��b"˫�3,�R��aq��5#�V��"DeZ����ZC�`$C+�})�'��,�<^���`Hb[�@����o{1oO!P��ED��5*��i������VJE���j"RZ!�4�Ñ\�wlcS$��;�ʱ�"Ai'�R�c��ЈC�bΗ9�4�!��91R~kC�@���`1�������aV���v�	`<��,f���T���3kl�`�t�r�K!9��t$ �
��2�";�Rg!���#@E΄�5� ���!I����I*(#�	��8J���`����i���z��T�m0�2+���q����bs�W�����2��:Cx�����/6^�@O�h��ԫ�*%��3g�DkP CvH�1:��2K�(�|��r����5�4� �HV!U���pv��%g~�0��ЪX�"[	w�c?��LB�򁡁�ұ.�m߾t|WDF�/r�*�0F�K77?�3E2;&Ӌ�n5p��#d`%Vb��Xoq	&q�`��m�U�f3�)"�@E�pA��j�Fe<���5dnJMu(
���GD��ȣJ��,�rK�h�I����"���ް�&�&%^����A9eS�p�Ɗp-0��ܔi�D�K ��;"bAx���R����ք4!�%�	$�W�*@��X��g�+w�$��v�
j#�nF�L(�җa3�ಹ�;�3P�]&� �M��*�'I�6o�(�C ��ߤ�<^c@��e����,�D�fqm�I~�"j\Q����1���'C:PF,�7j{i��!8���1�ma��6��sZ�2�����h�-�x��֠�d7��;.�d,�L�F��P��D���zѰ�;`���M��Y��4�ؒ��Z�F�hc#$��uˢXZ�df�i���4�Ё�&k9�nwƐP�$w�L�ӼC&	*~z$%��3W2#��&�MĪ��Z�4�a�QA�!���ڑ� ���f1�gM ��"�1�-�кyܓnƣN!($���~HX�l���CC�"ۚ���A!؜Mc�7!#0&�v��̑�$� ��?C��p��Iǐ� ���Q�N��RX�!�v}�<�Zr�~����v��.���F����Ǖ��K�%�/x��M�E#�^�fNDFSe�
�����^%��Pfj ��g��oA����9���M�`R�I�:A��k2Dw��u8TT �,��l��К@7�[�4�q_I���4��[���3peГeBWL��.Xh[�����ߗU .�r^x�9� �&�^sn~� Q<���Fm��ќb��L���K��� pD�i4�a�Y��Vx���y�#=x���y��O�v��_M��MM�ß�T�i����bB^I�'��4� g	{�Muѐ��;c{�\�˦���XΞ��dUbg��fM�`8�8��.�#:9���r���W�BmS�����)�aB@CrPnA����p!�b��B�̕�a�η�0�����P�J��F^�.���I����"��js[�"�V-�.2� .7b�"��� ̋^��W�A���8v����#�P�D���ԹQ[�+�7�FdX���c>�d�� w�8�\:�T�bj9c�zΞ��r��,a�G8�� uw�������u]����2�3�N(�઎Y@L��Β���V�r\��^��J��m#��wb@]��f!㼠Q$6hU.ó�
�P�l�P��>��X�hQ�G���Q�2�z�ӡ��(�FJ�4k����u鈴v��1���2�/@	2�Jf5;�7O�:�h��a��������"&9��J�@���#�p��C$�cj�jZњ���MĨ���<YE�u�(Nf?��S<��t�@�Uʽ�����'�q8U>���;�� -B�Q�.ϩ�m�"�����W��M5�����72fFZ��j�
�M��;'MD7�eRͿ�F"%�d����(��<�gA/ 
 �d��Ntx��(m�Q��  ��U��Pb��)R�@�B��H
�b��[������A�f�uZAM�0S�y�w�i�X/�v���B*=d�����i@ܾ��� I+�w��/KDg(���զ]"Rx�2"I �x�]*	�bk�x���!�p,�;i��ۉ��4JO��΍�'6� z���ѕ�c���3���15����΄������Ƣ2r���d@����FX�F\�9�K�R�EI��ЉL�W�`���|�H�!����JTd�{U�t`�}3��bnN��0yL2Q���@�`bP ���v"4��Ԙ���4��-!��3��I�G	�bR�<NX%G1$�Ɠ�	 ���HH'�,R&a���*��H�U�͐?y�=-�Z��!F&G7�"q(rS��t�`ܰZENK��Ƥ/%� ��?&�8*�&}6�ԍ3;�А�7�l����V=~�? �I���c� ��M�l^*�EW0��K2��cP�!@�l�$*�F�T	��/���(�b#�7�xH){L�/Fx�hr�
 q�W�dJ����V�%X3����&MO����y�:q�Ȉw⤹환��``�s��5;,�&1�fdJ��g��l�i%b�_�Z����/:2)e�ϕ�3�΂�{�m^�ޢg�@		`��;g����irL��Ө�!d��̝\.��E�
:_�����Q��}���1��m� *Fl�����2K����j�e�7'D��Ea�1gߘh�����X߹}Y��L2%2�!¥tA��D6H��j�D.0����	L���7g��=42�ۓ=3>3��`�hzV��t+��@1�Z��H�a��Z�h{�+;��~{� *=��ύIJ��h����j@Q��5+꿈�v��Wk�@"��"��=�� $#(�k�{�z�$���CR�b�̉���{AUd��C�����FdY�l9��9��Fz�{�YC�IY�z4�+2,�1�h�K��� �q1x�:V�s+j�;�4�c��;�駑(����ܟ��`2�KW���Y
�1+$Li'�B���%��hL�)�c@�.�j�F&� ���2�^+�fw�M
�P"�@����Yq@G?��ؕT!
�"^4.pj6}�=��P�B�e�vn	ۙ��t�O�w?�i� �/����B�K$Y�>�?�I`���cVt���j���H�1h
UQ�$6�4�H��ngX�r�p�����ǟ�:�`z/�H
�e�?/Q DGt�oi��.����~��f C��l�Ф�
PP����&	�+��N2i4�/�7+8𢡄OGs�ߞ^4 �7y秗J����8���j|z�`E�T�#�4Ua��[���K�&i�>e�5apH�`I��tBb K=+&�1��A�1i6�o:(���UU2L��� bG�_Z���H���H?�Zo,_H�DAkZV�Cm�Cw�
�C#*v���"��i$�L�m#��$�0 u�q��a��  q11R��!B	�*d��3RXJAH6I552Q �J�0��| ���Hb�'Y�JMʕir��E*�=��k�@��A0)d�U��
DL��Ă
]�(<*`
܀&K	H��#����  $���\��ƋB@��cit�������F�f�����߂� 72���[�Na,J������(Ā+m̌-�u�2����*h�g@6�@FXE\ĥ�M�M���(��i#��G�G��)��zgK}.>e�o"J4DQ����V"p"�����l����f7�v�^���;�<_;��Ҿ�,���I��6S�3�V�ф,����ڽ:�Y�}'�p�����ңN�E�t��F�ձ�:�CRXn|�.z�В\�&eb�	��AP�������PRS>���-�0l�%�*B--���95A��Fv,K�1�)	�b"��� zU�` 0 �a1�kS�:Vj7��'�&EIH�ͼ��r�0�!��s]L���%nLf;���7*�$V���aΉ����@��V$	�S�>��0�Al�t;s)����i��&w;1m����x3�$I(��Ȝ�� J�]�<w��D]��b$�Ɖ̈��{�u��	-H
�,��20&p[��ꥨ�(�A���FO9�W�,� D��xq�.�&@"90���2\b�����t7:Z ��2��s{oz5B��L����YX�& b�dr4���� 7Ā��!HR�
ɡ�N]FS�M �u8V2"ѽ1Ͼ����-:�� ��\p�
���v��� ;�v'7�6���B$�DԎ�.@�	J]�f
ԁ�ReF����%�ژs���*[����}�j#��i���ĥ��FbR�$���JF��ܮ���Hz�L\v��y�IP�$!��^����Y�0��(R@����l}�e$"�ڞO;�e\�\-תzjrX�x'1;��a�$��)��[o�:�۲pց�1<����+�SН��kT�5Ԟ+�b�@u禡�̺�+��63b� r�2 �u8�4[����k �3��?��f�ȍ�:�C���\7Dh��6��3��ƉR�d� ���t��E�2���NK fa�J*�c�2�g�'��kJ��,����ЩD��b���H�<���"xF+ ��J�����Sɜ	������r�2Fg6�|�`D9Ȇej9�����@�yã��7�&I�[�B��G>{-ћ�(0"!�eF׎Dg�`���$Ɨ�1 ��pQ���Т�,� S5�A�)��<�#Vr+@d��N��!U��*�vt0-,�܎"A�,�%sr�]Â�H�EC����D��f%-"f4�90��T�{jP�@�
�����MB�����d��ƥ4� o�&l�Zj��0��;����D11���834h֝��O5.����Э*DBH���QZ$��a��!*���&J���@����ʵ_m��1���΅�	���3 �Hp���؝����49�K���@dN�߆08J���g�����&we"=\E�fHa����N��d@�W���u��u �1�\|%hA���y��k=�*�9�C��kXt�+�{u�:�4�"� �[��gT��}3S��m9s�I��[�N�!f����13	Q����բZ���N:#��3��R 
�-?���T,�O}���r�!�k��P@Ҋ����M��AH
Dbv�g��B�p�C���M6����#;��7H	��מbt�06�۝���Dk8�a�$4v^&j|� �N#[��bUHA��F5�\�c��ܦ�8@-����z��J �o.�L��ּ�/J"�;�j؃#h���#C��ELIyy�X"�&����iL �t9|pN��H��Y�c�Md���9�:X ���B�lA�HO���[;ބ!$CF[=[�B��L��2����"Ȼ��*t��'��O;���)��ӬLV43,�2����~���X�/��]o�.C%{�g9�:5rw{��x��Xƛ�uH{^�0�z������+�צ��Y���*�gj��1H(ܨcm���E�,���!VG¥���� Ob�L��Aϣ��	u'"�����&�f������ldb����zLJ0JY������ȁ���^�� �����d�ϙtIG$�/��ޠR	!��ݽ!9�� ##��C9�t ��(���8�0��L�H�Ǘ�b�z�m:�9 �7'��ܭ%�Qp�w��ƙĖH=��w�ꡅY��?���H�F�ē�\������� b�w�׍ T��aI�$�)@`K6�n{��	]{��o�s7S��Kz'ͳ��( �ۮcV�2����ꃛ8����<���I�,�u#����ѷz�����A��:U����m�Y�L#�lv�;Ͼ���O�CR��F9O��u+�~��1_ޖ���(� x��ח��F��>���+?XVm��Gm4@�,t�ϗF��2�U��韜hT�{�d��@s7>�=1�0��|�������Nq��TPv��{=� ���;<:� �S��@3�+�B���a����Q3���-�ƣ@a�f96㾫�"���}� �'?�#� ������
 ��:s@-��mr�iG��m���5L�iŖ�'��䡖&�� U1�^����y��:��C�q���;A�0�E:�vcՏ�������|�i	,��g�������I�!p.�>|���&H�����'��~5Z '�����?=:�&yOOc�+/@��@�m�6#�Q ��c�<��Vw������O�3�K�z�y�&���ŵ�e7Ͽ��F�J_G)c��Y:K.�z˞^����T�����m/�'/o�D�To����e�k������Е�Z�x��1qz"X��Ì_=��J�Q"�3yX�I�$�D��cN�ʉ�I����H�DM�63_M
��@DLS��K�&R�8���q���g3W6�j�E�����ư�B�x���N�u���P�Cx	��q�1x�  ��O��HTOh�5�J�>8Ǧ�*��G��@0|���{w���գ���ΠELc,z��F��� <��Ύgw�D(���Dʐ����ƁZLC��7��uU'�l����1Sgc�ʹ��=_��ao��A,{�*"s���%�Q���S����FD�υ��i(NF�k��I���t�Z$�)�� ��Ɔ��B�2�&8�HN2��e��9˪�.@�0�E$�Z@3�=;ǉz}% �����V�9�q�Y ��N�t�4��aNw��ύd��.��+t�����f�=&��7��c3�"x�6��LD�����MA 2,7�q�ƒ���%0s;y���O����B�1n'�t�V���%��j���D�mOݍ-��'��#��t��y���:�]��m�rS'NDpLf�ȃ�� :?x�z&+>}�:t�eҿ��tጏ���.d5(� �S�-���QȠ�ر9�1�K{��&q��Yw��~� :8A�K��>ѭ�>�u71y���A����j�CHe>� m=����X c?��s��Qm?83��Q0�>[�>]U[�|���o��h-��ϛh@�o�?Ӻ�`Y��N^�oN�x'����0�v�؍�$�'��dH�$Bgh��(�P6UbK��Ʒ�Fw�^��],�I2��+=Σ�3��up��n!d2A+��ƣ�|��A ��'|:P��f���mK0�S��B:3��"OD���V�b�T���ce3�ovw �@��pn��[<�?�S9с&n�<m�-�EՓޥٓDX�h&L ����сL)��/0���2��e�N���H�vX���;��ʻMv�� �����Fԟ���Ma)����k�u-��I�x��취ȊIBN��G5��8$��m��=	�R=,����[I�"�9�ҷ8 n��[ͬo�����.�1Sczhܼ��=37Αl���Ǥ�qlh�8�V6��v�<�'%�;��xq�`��@�	����iC/M'kҸR��c	�Ʀ�/3ﮬT��`�+Io=��=_޽'�g�/���U��/:^ C���������qz����P��?3�D�`��^� ӛ�'�Ȼ:�e�BI$TF�Y:�#��@u3�0dK|���m�욃�r���"����D�� �\��0���nNH���L  P��I� ��B؀����‘�NNL�]P�m$jBČh��pJ7�4\�s���4L���lgK��9�eY16l��*Ϙ�+6�#81�6���\ָ��0�O3��H��!��<x�Հ�`���1�� �k$�� 	$[;_=�w�p'pC��%&3,Lvu3=b��JV1;佸�M!
\q�\L�^�7(c$1п���B
f��n�:�!h,�(�o;�5"�6��[�񦍐y||�u��b{ǎ�a2a�����p���'�8�%,��z/��P$��6�<i"&vЬ�n9���Z�ޡ��i8��������K����֦��{�Σ�P����^��D�/��#��'��1_Z����]'h����) ^�J)Ӯ�~�ۯޡ;��ފ�=�J�i�]D���E�4U(��h�qZ�fY��s��@NqD�:Kzq�II2�ڢ�aJe6�i[G�i(���"TŒ�i"��20�l�Ð/P����Wq �'��;�QBò���h���H���D8��� bO�N�Pg
�"%���<��	"r'���%��`~m� � +o�C�a����هHH�fw8�����@ba`��}�&4B)<���/�B�zf{t�]%i(r0I�+y�ep��ϓޫL&��XE�K�8u��L 32��0��J������R��}��*h��m���Ɗ�N�d�Ѿ���KeB#�|}�J���"��8��mD;�P�z���!���x�N�UǏ?6�S`���/V�����F��������H74���54���x��Ʀ��tg��]P���Ψ�>Ew�� 
������S����^]*�g3�%��Z��
JL�h�m�h�)$�� e��%�ўLB����hL�*F���*��=	I	P�����	� ��J�Aw�UY�p�'&2J��\P8�A��,�I�P��	�: �*�sS��A%�� ��n�
	��{��'�e�z��x��U���w%�^j�"�q�vlcP\0���/�s���ڝn1TLEI�}v'8Y�)��R#(;c�s_�$&8q�Y�O�$T�K�����N�@���x�%ff��tL���ZS)��NA�^t�l TdOi���􌉲�;����[�9����L�Iam��x�Wt�LZ���fM�\�8���)�1��zGVrݭ���7.� H"0�]���ԅHt�H�m�����5~/�M��MA����A���/��Ǳ��I����!����ɝ@�J�o��0)��VID �I��7|р�<A��:u�|��h���`���z���Z�2\���L"��J�|FHƧC*���4�67Ѣ �#(T+	��MIPYI�����D�%')��:�$�T���Nt�1�o���;w @7�� S�2��'�po���R�g��� �j�f;����I�X����hվ)+�t`KL�+��Q�%�G��/�9� Td��Ђ���c�:@J�j��o��ш�tD�)�z_�	�����QY����?$P��e�Hݫ�������gͧI,�=ѳ}�wH��&	�.�1i9%p��Z�|ZzTo����wҿ��+w��o�e)�y��T�fy��^�p"L>�ݍ1J���Q�<�<Ƨ����1׶��b����vϷ�'��'���h9���?z��0|���Ӕy�Z���������ND��y[t�Ԗ�M�w=G!�L �_�o��XKr5��5:l� ��sW��E�
:ќ�煉�wڷ���}�PD̯�>����9̾5D2�Mz]4�d�W�)��x��;����Sd��^ڙS ��״u�$�l��Բޚ�~�D� �[A�����������b�D���6��rN�\�ڒ5c/���Ƥ"��꒖��&0y����;ϝ		 �'$^�L�6 ��<Ƃ��H!"�G]��M�!���CY7D��W��ڴZG��ѿi�2�p c2�����wi����g�x�,�@đ8�~�M�12~�x��'�}v�t���iO9��{�������6���p��||��Aà������fU\�~�Ǎ��z��ƺK��<�  � ��?�H���%�o;��(�롋5r^{21�Ɯ;�1;|�T�Z�S�0L�m��%�v��H�^+����b������o���T�=� (�F`g՘�H[N���� @�M*\I$n<G���X掟+P�$����c��?:�K>�;tт�oW�3����IF����4�pa��0yVt*"�Bq1P������v�(��8}?_X����X�?���� ����	\����i�{��jd0D����MR��UҬ}D$G���G;jv�08��ͱ�М �!7gs�qL�Q2�U\d|Gra&y���mL�e����~����c���gB$�{�u���dgz������5��xb\�].���,1��L����n�XgBq"f��r�{�4��#�O!```34"�6�4"D#Ib<���j<@��O�|�4$���>��H��}#x��P��Iw3�e>|���t�J�$�6Ԏ��_X���AHw1�t�bm���C"F2���:\�eB�g,&�2-�8���������x�W;��f�t�tPa�\�;��H ��x�Wa m�@�9�7:����MΙ(��E��MZ�D��۱��<T�`f$� �3�t<]@���Jf$�D�`���X �N.J
�ı)@�����M��/K��\(@9&�O�Up@��f5�:��C6`�Rj�F�Y��k1�)��'`�� �R$����S���K�q���2�-vǼh0TRGi�	q�/�f�W}/'.��j�=kOh&bSi��L��T�Ȧ6E�G6)e���DS7Y�9�V ��;�;^�� H+!�qY[��@���t`N���1�ؘ�`<I�4:���FSvJ�P19�e��h(��Z\l�0-� &��Lb��2L��K�[!�rM��g!2ۈ#@̸vJ<�cX�(�
�3���BK<��M)p�5�	�z��N/���ʝ���:�8JjԎ��a^�7��0�ӿ��jV<�g缟U��,3�E,v?�����&z��_�������$$G�L$�3��w��W��ϥ�.m���c4�q��vZ��?Z��X�n�6�ӗ�U��X����"��aQs��$�ŲLTRab8�� @\�R�1�Nc|a)9L�n#�\r� ��9���ɤ�BA]Fc�c#	̒[m�"�g2�(�:/Vf*�"�+��΀�%�v.�ͣP��`��vv���mIک��ɩ�h���X�$��HV
���5�1�ED@�:��Jz�Uw	&h�jtЍ�b�%!� �Um� ,a��� �KU��x�d��� G�-҈�^�!�;i4�r�1�[T�'aA�!��`X�����T��H. &zkq�'
BPótA�P�%M���:�d���P�ȫ �Q�}7�Y��U߼�bo�9�zV��+ ��&����%2���1L��7�u�}��jc��ΐJ�fj}��]gA�����I��S񝵙�&K'l���� ���j�]��5'dU�_�+}��;�̑E�<��5�5���#��C�8�qI� ٬L�4�����r����y9e��� �;�1{^��I�V��/C��)����S��:V�0K�4ț�l �&R5�$�-T�P�D!�s�'k�]N��jK�h�B3lN6�Bd�(��d�Y�vK�SbKDZ�
e&9A0ɞ�"�K`��DhC� �B�c�Kp  ������x�� l�(��c4YNE�P�@1l�~b<h������X 4�}(f!R��8��\�H	� �� $V\����C��B�I*�Sk"җ�CIFo@��	�a�*t�#va%�("�V�M�Y;���F8���n���2+��"!4j ��wf�4�*���b����B�{�s�i���rgR�%q�RC��,��9�v�OGL�
Kc��-E��3uo�F#
�kG�b��������"7#���s�(��ð�0�Rd��[�)���ci4Q�5�ǳ�h3 ;���h�l�:�l"<��D�J���<�E�:� S����8�b~����O	�,U�ߴh`6��q[�5ك�_�� ���eH��+��ER'�ܬc�Ja1�JL�zx�$�6` �,�������qz=��$ �3+} ����M�$Hw�h}YG@00��*���� �LŅ֙��ب�!@JF�[��&d�P�2�d����7[���	Q�mh�8	�+��3����/�d ���Jդ��k$�l�T�4��b�5s��"R� �H�5%޳�@%�W�Y�ruF#��ሂ�q�VH��':�(sq�(�Y�"�� �F+�Ƨ�0L7�!G:x���fQ�r!�ԍR" ����12�:�@K�z���ٓ�Ar)�Q�B�@��ͣf �� �)Qdb$1�x�I��I�쁩���bq2g��0F
]sX�`Cc�%���V˵���BIN�i���`�`kJ8 ba��zu�Q�b�!�Mp}A^�-5	�`ĳ����N&�f�k���1s�W��`��j��i��N���&:��Qf#�mY@��sף�3s�>�禁VC\��1���I�Y��^��DiW/ϟ(�HP�h��#�G�qۣ�
F�y���WpQ,�l%���&�.RL�(����y��H,f�b�K=�ny1GA�kD�e8�[9F��jD����R��R�a$@""�d�Zפt�li�޲�Lm8�c�4q��.�-�Z$�*�¿�LMV�u�T��b�R�)��		BV'���F�@ ��*��� _4r�M��E� "fX
�GL��e|�[�fB��q[����ٙ�7�0��`��*0�EF�Pk�C ��#�kR��0HA�;�[�@A�db�ع�B,��
�o	���f&��p�F�8��E���.�1��}1ڵx-�"�Yfm͚����C'<�H�j8������-q�V҆7��
32.o��L/��A��� �C"�]�l�F�Ab�W:
�
�`  �h@��.+%r���Ĩe��߶��iYv�g��jA�u���k��)$��"Yn�mEEH�#7���n�� V���}���!N�ȏ� �a��%��ôw�J2�I����n��q1����Þ� B�$�|oET���_$E�V�㏾�1M�]q�K`�lv?����d"#���!q �<�b%��A{It{)$ �m��VT`Fxa�	�.m���A�B�44S0<mff�m���ʢ�����`K���uIY�%$I��qh��(]�"� ,�Lp���F�i�I%#QM��E�-��@��#4�,�B2�6��p:P�x		9�6F,=�a
��eF�����n\08[��]j��Q�$eu �3b��u<�j	PJ����L� ���D�D�i���pĊ�X�S&�8(�+A�0����.4� p2�M�cѸљ�v��G�>R�\őg��*R�m8����Թ$x� ��ھ����+�q~ �f�p����{�DJ���XR#����b���I�B�O��S6W��zy΂�>������5v�5 Ҙ$�$E�F���d�KXw���%eC��u 1Ő�D�j�&��������%o 4NU���i�t&@Q ��9�AIDDT�K�a%�"�B�IP�V���}����̂U89H�`�iPk�c%F;�n4�thX�	R@���6Һ �eWQ�^ȢD����a+��1�m�`T֎F<���$��S�GS$L�o�����S_>�A��ӍB������JΣ
X�U�f�JX����KI���#ƶL���9��I�t�������s�1|:s�3p�(BB���gT�4� -�C��1�Lxi� Ě�J�5
 ��VY��������gP���d$h�Q�A�� #=�l( �
�$���Γv1�0ƍ�#2�.I�UfeN����$�MC�QIbI�8� �Vlc�n35
�I�Z�>LI
@��� �f��
cnB���q���UBm9U�!,�>#�^�l�� Lt�TV4A�D�1G'���ϟmH���ҳ�m,�*GH���:t��fb]�O�S.W��V>u H����'L�d�lnn7?ޣ�1\����WǄ�8Q��v+�m@�RD$����P %%5���*�X
D��}T��-�d���Ӈ�@�2$��'h�0�H�2��0-P2�&'hE �@�R�Yo�Fł� ��ݝ%=�D� ���CD�A��w��F�3DU;�7,�3��G��t�B��0Dh�d` DA ���L���� ��P���K�>�j`RB�,��c��I�2g�>~�(3M�e�~q����|�����Y��*��4a�jRW���Z�f`���1&�:��	J����jL����}�D��eҾN� ����s���J�e�"X��|V�uS�prI����>�³�ҳ�dJ�Xs���S|���ɶ����<��,�d��b�Q�/����vs��5$"���N����R@[�b$獹�f���f���\Hv~6�L4�둁U9z��]�A�<��H#l\I	V���#�1���n���:�d� [�mH+s�%[��wi��*qܙ63�\gN�@#��ϒ�cx�g��,K���l�)9b]�1�L�@�9�����C�Ͼ�*T���3��t@���f���Y������j1BX��X� �ids���<�(��ܧX�=�J�b������A;����dCi8"g?{�9@a�a��,��V Y�(L�~�S�P��t�3�+(U�4=��DN������ϟ��<?8ԎX &	��|�ӊA(�^ݿQyws|�{�,��m)J���o]�'M* ������w �&��qM*�3�Й$��$I���&O$qJ�K(�<��YaŰXu��8
Dl��x�͠ab����A$ 	���<+��=�����A$D�L�#�А*f1�Ln}��Z�w���.���{���F$�A5eXl��ҏ,L��(�X(醔@,�O$PFWTt@� n3��0�P�����'��M[2�(N@�(�h��W��΢�b��+-gâ����BS��+",-M�����d�"���t�5u;����Q�m��/�;�%@F����e�i`��jg�D�ܛz|��@�iYbv�*v�y�D	��ji,�l?�P;�v���cfoNTX&���ZG,@J^m�!$��o`�7U<��cd_d��ȅ�s/Q !.p�z��D��U�����\� ��HHw�)��!	��Y9%��r�:�w8E�� �"i��E N�BrΆ�$1[	���@y($�L�Ew�i��������;������\�Q�������4�:4��^mH��� F ����lh&/1���Y���p��
��KD�%(01% �щ�8���
�C#��D�-,��&A��$�Y�bo}z��t�������F�o��HQR�����pq��(�?U}�{��ɏ�3�A,s�F�&Ҏ}��cq7	�JX��tm�$��-+�ՆNH�3�tP9K*#�}̺X���т��-���Ed(�H!�H��K�`:�`�
.A�d�s 2�� 0�0�"R&7��Ϥ�x�����+b��h�a�hE����wΗ99)���x$��^����TI�#�}M3�j	K�b���H� Hn�EJ�`T@����Z`�(oߝ�S0�RM$�Mʹ������DaN>�����'��d�y�r��x��z�ɠ�*�K� ��M�����2��	��!D?�dDJE��\!$�$RB��d%(�Vؔ˶�����r�-�h�rM�)A�a��
!�Mt6瞺����l��7��#H��<9�դ�z��v�#x�D#�q�ᘎ� �&�����D�O&�`T�1�H�V�`�$3Qw�t�WM3]jH����`�w߯M� �5�`'���}�بߝ��w�l�$E����:�ǧ"NF"��"3��D	�po��)�(��P�H��T( HC�r��1�7�2�GP���~�~H
�[�v^]9j/�H0�JX'�ILs �@�-�/��� %R�-��K� ,(��:��9JP�T`<J�#�4�^��f����E-6g��(Vz�vy�zL^��l��&!�ŹQ��!*�d���c���D`z���X\V��RZ����F��B&��#R�h��M�bő4��î	#����zjt�"9ly��i$CL&����K%'���|�!�Y�Lx��2T�����z@& %y���P.��7� 9�;���"��l3�W���Ւ��׹}�)%�o��<��P6K� �T ��x4����[�5���z�}*��dv�7ߤ�AyR(b�=�M0	�`����#U�0/�D	�!��E�s�1QEL'�X��5���<l�	�\CoGw�v*���H� �܄�|b&M�j_��
į*��cP�t�	ܽ:A�h��gS�s IJ�1�D� ������a�ru�_�@!S%�<�i��("w���ۣ��w��(�1�He��)�5Xh'�3�G2̙s�� ������^FFW!_�n�LUe�qzA�+��F�����Wrȓ35��� ��n�O�B[�ϜꙒ���>t���;��y���QE9�:rwRCH	�s}���a�"���΢���R{��\cRT�_����!��8,:A^��As�����B��<s�R)/�~X�h�* ��������8{���1��Λ���71Z� 9c���N�l�g���)5��� :����$+*e�~q�� � `�$v�gC�{"|�e�c���Ue���%���

��F���5VL v�� �à`d��؏֠B%��o�1֏�Va
��c��1�k�qT����U�g��m�u����<ߧ:�Vյo0��p�3�L�=Y�ݎ^}�@ ��� �	&�0{s� 5Aa�߱>�:Pe���ә�Q9������M��w�7��i�A�L�,�эav_55!$�H�Ќ�Fy���.�>s�}(���>�c�����K��Է�1?�hz`�_�C.��'����N��?>b���۷�^�y� �Ck��3�N�Ƃ�T��s�&��1=����g�����D�CpHɜA�*��bWc�b#D��4g��ˣ��g�c���@����p��I�8���bM��z�7�/@�"7��MO��͙1$^#~t�d�$e�X���m��b�T��	g<��5"�
."�����/�q�XMD�P����&`m����&.�N��gQ�w�ފ 	_m�f3��E79�ޗ3�X�z���za�-�A��=cI2 w"<�P�1��d����x~��&k@�7Lo��K4�03�{N����:�q.|eБ	�v����%'q��:�L�V��uԂLw������LT�+�驨�����.�ƭq��J�pE��)]�f����	T�Kv7��ߍ4�[������cƌ����_�G�e`��"�)[���HĲ�qޣ�B$�kx�3���d��ϟ7�NP>~]D0�L�k>�T���������R��88�e5k�"6�jB���7�Y_Y�ٛbh�<D�Ua2�-IT=Uo�a@ag5Omzؖ1�q��t��G;޶="b�n���W̷���$
^8n���9_!"%�����՛������ВG&l淆�'��B���cf�rs�P�J���8.�Af�j&6�T쉠���1�*2F=�������ӡ�-rf'�c} 1�e���e�4u2,U���t�0.�H�,L.W���;�<�Z;l�/��e���ML�X�LF��/�y�J��ً�&p5$<�,����0SPq��7�X�
	- /֣ɤ[�H#�1q�/RI��#����IЕ ���r���!2UR��U8��ר�/,��r"o�� ̚�#�����*�@01�z�RCa�j*��� s�,�UF
�wqҌT�a�\Q��vb*)Զ���sp�"�r���E.���1`�y]��� �L�c<Q��%��M�:o}�U帘v���̈́��Xb9;�ۙ�0���2Ff�{�� ̠F�*V��cK%#��	�B�&̍��"v���I�B��e9H���c/i>��Ər q�`��$��*N���j$	(�s��$,��4ĸ8�=���ތ�J��G�:E���D�Pb��ޔb�3s���C���J1~ڭ٠�.Y�y붪��.�8z�6X*��9��58V��6��\��2c+ǎ`�l�[IѼ���dBB���Db�v4b��Q���i�;�IX��d�(c
Dڤ�=+���&��N����W`
K�b��ά�#W<�|�%�I�3�75�!�c?{�E�������闼v��{i��l�="&�� ��<�X�ΐx����^��*����L7�z�[{n�fv�5�m�T�(�H!%j[y�۩���ˮx�=I�;%c��7�]Z�b����}P�X��nv�u�$X��3��PI�
D7i�]�f�>]�df�Da@hԲ�G9�QQI�3��t�qBI��!��4\%�#�$����/RP��n��S؂� ڧ��٥��Y���|LD�hr���Bf|���*xɱ㦕�b������kI��w�w�@�崶1� n;�\E`�&0Pk�s��6jPLq������	x��~������<m���33�ފW��%J���3�#B��.�-/�ՙВL�{,9龌U�V���"�H1���� ��-�4���EVz㾝%�M��s����N'�5�ңrI��x3�BڳJgFu	���강c�uq3��\%%NY�,�5��f���1>�(;޿� ,&�y���Y���/�MHȎ�%�|u!gX)����n��]������|�Ɔ��w�ݟM�H�����Ld
��X��Ր��{~k��1=���H"-�y��t�

XSy�g�UX	h���~�#Ʌ��w@B�n��W��F'��M�fL���wj�&�:Rf$]�x�lԠ�Py�Dݓ���t5�'(n�g�5@�˝�=޹��s&}c�#O!A¢+�}�H%�Yv;A.�0Dl%�D퉼Ʀ	f�_+��/L�m�b?�U����kK-�輾�;iFm�{w�h��Cn�FW��#C"�{�Ε5��;"#�/p��̚���	�fW�N��߶O̜ 0T�_��Y�Ae*�:^ci�pE�Z�n����-,ڀ�g�Z�Ѻ\�M�Mۨb�<q��e8��8�I����צ���i��汿�I$DU�t:~{}`�'�c���DA�H�K��X��&dmA�d`��>W� v-&ױ\8
"���G��q��u9�+���h(
]�<�<�W��ǟ��@0��ΐS�^�\�@(Vf������P�
�/�{�X���
���4��n��H�k`yy'��9��#�{�y���߳ҧ�H�V;�޻i�b�g��'v�U�r��$ț����� �D�p����ćz˷�SA,�o�M((0�U`���bD���<����C9��!��~��Pc�Ng�gM�ji3��w�,
�ƍ�����}�.rQݛ��ȉc2M�!�ZX`^����j�(akM�E}�P���55�}w���	�ٙm�V,���8��ٝ�L�Y�Px7�5��A0V
t��q��+a�������|����Q2�ɞ�yh�aTɠ���u�$ȜN��b��>��[t�b��ɹ�W6 �$E��	@^�/}�u���D�ca�o��s`'���aBl�p+0m[5|92�LE���\�r`S#�L��>��2���6i�Sq}�>C�Cw�J�}��@g$�w�l�r����Z��Ϸ�t$N��!�L���-V?���MAo[��(L�o�G�i�-��y�7ٽ
Dp��{�2e�_��t�t���Z���O���LBK-'i���Z9D⪎~o�$�� /���ꂉ�r�q�>@� ��X�{Q�BC;15�:��!���i��X��v����������{`)�=��"L�4��ƈ� �f���	����A�!������t�P�m��8+~��	��L�'g;]��:��`�7���z�P,G{}I`���d��&X��8��,�g�DK�_�F��HR 篮�`(��7c�����"HSz��%�N0Nd�s�s2���_�����=7���uRE7��m�,DY;sU��2���)�W��4 � q��Nc<�{��%a�۾�9	cu�)�Ј���\tkJ ��O$��ޓ���Ip��8�ө6�tw�?֣�o�~F��e�j����hpG�vx�tn�h �B�HәȖ6����t�a5�����Bl���[�,�~4�T����^�h" Z9���r�F����t��}���x�L�I6��s�HZew�ǜ�В	]��ϣ�;i���]���tuHK��OV��__���j��x
���
^��ky*d�bJ���v�8K,[�� �?�7�zJ�2���W7U��D�����:"RQ�L�@w�hxI�3^�2A�̴����rWm)��v��O���'��)�������}&$��JM�+��aΈ#�>g��S(�A��󞺖 �������������|�*����t�N��7�ƚ�M�ˆ�3#7��2�\3���&6���L��;h	a\����������gl���vm��Y�N�槜�.���D	k�Ƙ%{�߼|�8������s���:(�L�>v�?S�VV*9�������꾇T�r	a�R���t�n�3��~��t�i�x���AH1G5<�>�f4��m@L����U@�.%���\��N�EP|�cE�S����9:�iӧ��R&`3���_��	�:E�1��fa��ۮT��E�d�-z�M���zd� 4�Qbx�Noi�xч;���E��v�q:�J���2��S�M�L3Y��x�@/ft)�M1/��4��]���F�eQ.����P`$�ƁH*��܎������˳�}�Ff1 ��joq:6H&3d��o�u����bR\��N҇c3�&wo������&��V]�^.�������v�AƦ����]oF���@X�L���G��%�;O]=�����Yp;����VyгIdD�[�q�����!��卵����{L�LHS��$�ߟ���_s:�ffgo���QoH[�� ����� :�x�}����͹�H�߾��	K�3���D�����v�)fr�\F��М!@��~�	$!��ztѱ37��^�'HL׊�7��i�!~�=<^�1&�_?ߣY(g�\��hhf�����Ǝ�=3�8�b1��f
bz���#��<�^+�];@�yj]�DK
�:���q3�DD$�M������)�G$�=�Ƅ�܎�K�o�%��C�w�mI���G�(#����HD��^�C�DO�1�453^~v�HIm����z;`A�����bg+io#���};QMMf�j;�	Y�'BH�Ι �`C_֜i�@;���<�g�d!���������h�qg�㞚k(K�<,����gH�#c/Y���jB@\���p�uTue�s3�+V�>/yy�2a�+ M\d�:�hbr�����䑳�bc��ۓ�Q-�V\Ǿ;uu<LWJo��յ$�%iAW��&�F>z��I����(D��s������x���} �M���^���(Q(��nڐQ�4���d��_:p|�+Ro���6��Tb����MXb9�ϊ���S^����ƌ�r �I�A�5T}N(�⾕����Ɵ�}�]�x�����������u㿏�T�F9�� �EIu�<�_����Y��{�d@WMω��L�#Dn��@^R.ӎ���B�&:%6������S�Y��=,��I�w�u.&��BS(�P�?z4�'6�g��,���y��dL�L�U4^��]8�J����p����� �̓�p���A��qY��I)���r4��Ѐ�!\,+?{+�R$"�?>��pe��>d�ު�n���|�O"�Caw;Y뾙H�YW)�I�kL�"��y�ڊ�
�J�D��ω����:P[;�r)��o�h �1��tj�5�����^�t$��`	������G;3-�F��!}F,�Y溣���u��G�����Ӫ��o���:���h	�`����^z���<�� u��8���{�����Ǭ��v,��Ts�co�$�\��ۧ�D�[�F)�W����%��5�Nw������Y�M0`�]�¼5��s�~�� @�{��}���u��j7��۝�5�������Lsr������0��c���y/�*��6
H���=ur�}��K!@B[@m�:��b���|�h{�C<N�t�&"t�y�[=��Xo��� IIĿm Q1�i���üL�֨MVyy���,	���e�Z��^Q�v�xf��.\��%�T��>�$%���q� �lv7l�
�K8��d�M��ƚB�lx�}#|t������]�H�%!�?=d�
�D.�:�dݡ9vWڴ��0��Ò1�� /�_�f�K�J�I�n>��Ť$dhs7�҉�0��r#1�H�R���q��'@
gnH�) ar���0��7#q�+hJ�Y�����Rc�"sS��BTMJcm�{8��%����{w�,�޼O�����Yabaw�gm�ϝC�϶��D����O���2U����y����� ��U�s��Ѳ�>I�|�&1�h���Gh��}�w�?D		�=|Iϋ҉ ��n��ƣl[n{cΚVb�f")���a;����z��ȴ��F\}@Q�V1�]�i~�L�k=հH�,���y�Q�.��S2Np]臂 �f��ΓJ'y6<�&�:D��B�e%�Ļ�Ƅ��6h�/���Ej��'�ƭ�b2�Y�cd3��^°J���V�͋��M~-Cd�9j�'�4
�I`:�]G���6,j�K:�#��b�^q��Q�E̍�\u͍vP����7�(ƒ)�l��˿H4�j�8C��ܘ�'����������se�ٛΨT�ȇ;H�x�"�	�w2s;Z4&���n9��ab'�ft��#m\9��ƋKNe�.Rm�&49 U��9'��)����n��t�ʨ��8�<��6�P
�̓듞ph ���r]�;�v�)�..V�|�r
��d���F�dB"� ��h�8](<��i�޳먫_5������#�v� �|�A!�N��|�3�o��ТUZf��.(��k!X�M4�c)�i/"�U��� F�~cx�%�S�.k"�la0(4P H@��uHUi"$�&�>���M�B��*D�V��@n��Si��̔��'����8б�EB��)�&�8��'R	�d�Θ���T��N��#Hͺ�	4�S?#l%��H.��rRȲn�a25��2��D�s"0�g�`�g��Y���`++�g"D�Z�e:-�{jN�>	"0&�˷/  ����1��\�b+�FI�a�brB5�4$I�C3
y�Z���8�$�ɡD� J��q���Tzq�&cKB ��o:��}��H�m�bx��5ajfg���T!�u��V�!D2�D��m����\�5j g|J�du�"5]d�q;t�v�����_z�g:&F�hB>y��{���^�T	3����9K�h폑����c�禓(��D������N��|��烊ދN�j���0@������,�L�R���[��B���P�O.g�i�p����%GN�Ɩ1��~���%���=e�5P��ŝ3�%ZqЪ���܄��4��gA����f�9��iզAP�j� mt��(�ى�b��D����7!���$@F=�6�cMBFeDY'�MDEP��`n9�Sb� .��h�Ԑ�`JXJ�H\�\�u� ��w�D4���4nFb�ІER�"���le&l��[���� x� =���Lm/]+�Q1;���C�"
�s�����ё��������̐a��Z�ӮD��wj~ђu ��?�ƅ�_�?9Ɩę��Ɨ�i���ߍ���G�Eđ0�N{hei0'7˓�@0��3�:�C
dL�D��4 ��Y2*��3.��Q���W6隬��|�^>�����GO��������h�����欦ʷ�V8�.X�~Y�h��տwB�����$NHՒ��B0�Ebt
p�$f��:D )C*�����_^�����o�HP�	��@�J��h��=���C"�����X������
@IR˜�4k �6��,l.��*Ů���U	PN��Z*��Y�ot�g�k���ؘ�3�wI!R��O]>x �兛t髉LZق7+Lxf�	��;F~����u�����q�
씗�	o�t���L Fd&��y�����N�=9s�>�BVgm��9���� �(�� \��q��{t�'fXr^��jt�
-�E�,L�6��h�+051�:Pr�	q��]S'���j=y�3]��u0s"Fj0�/B�7��Q.S����ê�S���qy�Ʋ1���s���8PB�6����Ґ
�Ro=����N!�����4Ҝ�N~�U\���K���~zj�_7�[38��!L��Ll�����B�dL�����}^A���Y߮�0��$��)
gAdHgp
��>tjH�la���&�*k��R;Y��&҉���w�03
;�o}C��AI0b#u� �P�(����zk���`&$B��4� p�ߘߜC��11V<�}�9��U�k���r$Jz�n믶�����9c� �����Ѹ�N���a��n�yt��,�����XUvF��Ϧ��l2��4���?�W�t�˞���I1	�>sƣJ��q����R��]mPG�EJ�WD/a�j��,,S�ύ��!'
�OH�i -�<]��}
�"`Pa��a�5L��K�q��!m����F6h�LI�����1�n5#���q� ���*3�1�ޏ}��)Cc���˫蜕�n��bx����.�h`<� .�GgH���>�P��^7�i�+�~U�y��2�'����h�m�����o�7�siљu�������Z5� �\�-^q:*Z�YbHf�!8��ň�U�����-3��R�A�������/��,�H
�&8�Xi�^B/�׋�b[$)O��3��"������-� ͢��T��cN@�"�$�[��IU�J��v�g�e�Fo7}�헛ѓ��Ba1u>o��IiS/��_:P 	
I�6�5a��&yq�QR�PD�MU%���o��*�C������w�#����\֐�ADO��,j`
0�{�2|� Yi-gl>��d$D�&`���Q�m���h}X%|�j�����6������G��(݀�i
���"���%���5_Ā�#dV�ܼ� �1��Qޯx]"�Q�GI�2a0���Z���h͛��h�c���f�`�
��|��	L�D{Y̺��t�u�^�%�����Bp�c��J�-Vӵ����DqЂq�K��0���,%��2'�U�&U(=~z��
����$��w뢻D���_h�h%[)��{0V$�ڂq��
J�g�X���9�XE**A����̤�<��|�l	���7��.�BlZowޜis}'xߖu0B@Hc�Q�i�0��cA~^�A)cb^c&�ڢ� Oߍ㯍$����	ߒ������,M�L�΢8zwL�$��|�c:
r3�X�N��� ]�j�;t-�B,����s֮P��J�H�v`vң�'X������1��p� R"\p��؈�.���U�7�<?�30����\�&����s�H"f�8���cP��e"�7(�ˤ���n�`�qF�&i(w ��ilِV�T�a�50�m��O�:`@vLt�흽(�D���vK�J�
���,{�Df�l �i��:��.E���P���� +��:(��&�p]gH��Tj�L�. �BY���n��t��Ҙ�$"�jbk�wB�3Iq�o3�K�S���g�e�b�or}|i:*Q�D�Nt��3<�u���N���7�#�֦M�K1��-�+?2�P X,A7�:��9�OLq렡3���I[��3:=;H�ܛ�;j##v���s�o�	r��~�li���h�{1W�j�����gB� ��DR�n�� ��3��#!іj�Ye���pF2�M�w�4�B�.��t��kX')�"w�`��$v���CtQ0d�=�46f�0�zc�r�ĠXf�j�2�6o̞��It۳�9�#F|n���ׇE\����L�:�0�(@��eo�q��� J@���}�x���"��1\v��`̢�b�YZ6��$@͒f2�#h�]IA�dSվ�EFVD-� 
晍%G(N3+�D��z�{��:t�G�bĕ�Z�8�c7J	M
.Z�3��E�+�����/N��Eln���qz\N0�����ZVȔJ�@��O
6B)�yoM���L+.w۾�j��.W��QiH�`�3�`ǈ�5��6��8�6�(%0��!A���"@�fz�2N5
��'"�E(s#e��I���e��j?����s�BN`���_|||�.����3���&�S2C><W�����U���:����/�3Z'C�78�^��  @k�]o|o{�wqs����OW����} s���$�%�nc��F��A�湌��}�M5�(bb�g�����+R6���tY�����t�n�����P�ŠJ�e8�0s-W��N�`���,�3�/I	�'&��箙� V�nad���0�!P�H5��zfqImp��@�I����,��[ZZ����UIsPL���t�s"#x��f�&0��("	�e�%�@�'��ˢ3�$B&H� iI7���� d����F�a�!'$[	�8�A�3��ڂ6�� �O,0��S�zQ��ϿCIUE�*#|���S7�ދYf�bt��I�!z1;Ɖ*�j��ڶ`5X���H&�NQ����;cA�rXDWm�F�DV���U�j��2�fދ���5� A���@���[On�@�OO�zν~q��?�@`���������M� ���O���Ē��n�t�Y��H6� -��yR�H�N�i	���g= t��-��bm�#�e��M �)�Ƃ8�o[����� ����}Ul �I2�����آg�g��@�eFcx�g:��Pv��x͵Π'2�E�e�N��L
BY�Ӟ�����<5Ey��68G��=�A)�7﫥�Cs����18$��.���pa Tr��r��Եo�_}�A-�Ǿ�D�7t��t� bK��('��KBhU���.�YHJ%�1��>�8 "e=�7��-�B7�hե�
��LtƐ⋐�L>w���a ଑�o���'@d|��0-ڞ��R�Їb?[jP0DA����Ɗg�)3� )���Lra��u�"�Ps��!��Ԕ�e9���:  �cqvy:���E%"8�cs���"@.�ֆU���d�[�5��ZEu�Ɵ&d���2��s�a��3�V�K�ޔ���Hr���۩���Q*�����p��?;�=_�  �Jό�gL�v��?���'"P���V�f��� I��M������})ʻ[�2UE�|��4�w׿{���0�z��d��\�_���m��ޞ,P�Rǜ1z��\���� +   !1 AQaq��������� @0P`�� ?� �sΤA¾�g�?��.�@�-�GO?q� )��pNt�x�q��C����h��X1\�JI�/�M���� ���O���_� �A�_������ǝ )��;�G�C������h��rj�#���b�=?���y���U��p���P&d�f�����=4H1'�e�ԭ�Y�&�gm�󈧉��z���8��qQ� Q(>��6��L�Rm����m椺�� �B�coM�"R�bz^��}"8	=#�y� K� j=x��O�J'l=��a@r&�5"""<�b�N0=e����G�Ӊ��h
Ȟ���2$�ϐ+N�²爗9ߥYR�(]Zsw[^L���M�j����e�����:����Ɣ%C��I��A<�9괸��
`,��t��	Bg���u3\H���E�����
�pO��P��41��޵,��0R��ˠ�R)K*b3����l�Sy^�ɸP�ۍ"%t���.a�}ƮH#3�����@91����3ƕd�T�\c��X�Qq~���/�����;J���	�m�z�J=(�2D�1�ޕTSb�8��`�)c�:I :��8�r�
bs�zhT�M��Ǎ㭩�A�!�z�iɣ��.��\�nSi���om&�����F���_�H�f�c���Z�#�\����lgFCu��c:XLHJ��ܸ"}t@���8먹��9�Y�ϥ�k" ���W8g���0�}�wy����]�t�Ǝ�!� ��	�&��B�	��FS���|�cd4�Q]FT��E ��a�c��d"$�z&P8	K2��P��e��elW�&�``��2McH��Ԃ��j�z�:�,�LCCn��`�*��s�q]2�$��=����U�w]K��nپc~q�0\3��s)�P@�F[.��N���N�S�6�57�i��1׳� ���È^s���iF� ������$��,!6�$���6�r0�h�h�3�Z4�`1��d�#�#b&��ƍ2pKR�8�Ơ���5�H��:�M5%%�d�m��d&.9i��W�D�g���gir�1(N��\C�uRn[w�uDb�Z^�q ,�Lmg]J�d;��\ n� ��,��D�n��K�a��x�Kp�T�*�U�#IС�HEl!�\ $A0^�g�iJ�RN��c��é����U�F]�HH#Lt3�,f�4*�wd��r�#ag�.�� ��[S�T	���
)�*\mΖU�Z�bx��JPXM&�a��chdBiSs��C8db]�Fm|�L!\($����]��kؠ���q;�iY�2hS {��#�sj$6n��T��]����ߘ|�3
T!��2c�	U�i����"� �fqz�QQ���x�z��#$i�7kmKy"2L-��C��R��̲�\&#vZU�D��2@���6�	�����V��Z~�eb<G�ۈ#FM�!��ЖD��^*$5mI#�::BB37Ojc�t6��w��Ǝ��JX�I-r��#"�Í�;�hJ��x�^�;��@D���Υvv�6��H�@�l����&�TN[�̢i�����}Gh^��b��''��L�x@�������\�#���gC��}�*�7���x!�1M����@p��K���4j*+-��}v�ӓ���/O֯`E�ɒ
�g<�֡(�;��G;@E��Yv�6�%s�أ����43�����DLC�#�\ɩD I�gJ�3d��2�Gn�@.�PAa��iD���D}qgv�6a�s��Ӷ�y-���� ΂]]i�6���65��7	�yҔ�0((8����4Lp�u�����a��~y�+y��,����LP��Ï�u�N�{_��T�jU�<��wv{DF'���H�������dR8��RnsN�Z8!",(�D����(,Il]^f6[���RR]���1$�o�;�*4>)��(�,:K��ɔ���Ɍ�E�v❠���=F���������$`A/1<��JT���,G/5�ҤQ���qe�tmP$�6R� ��:ÝBS����ӘV�K��{:p1�h���I2T�f�7��xѲ,������
s�)���t�jJ2M8H��4e<������i�@�/���٪� ����oww�$g����c�=4���a����ꡃ��y��0��==;;�H;�c�^9�S�GK-���"o�^�7��0l�ܳsƁ:3l��K���;��q�l��	`"�q2S��'��`HD�F�:��V9S�Zw�O�& ����x�(*�v2���芤�&`��#'}Y���b�MS�&�8�k���"��)U���E<[P�R��Vҝ�ץސ�$������p�$!#��\��NG
�����F8�=ȂMa|߀̷%P}�����-�:�}�{�.L�Sظ���P�)I���Ɛ`��`���3AP����֐�ҋ��AF�z3[>��o����s�3��,��x�xй���.i��}/S6�����M�j�Q�^A�D��ܝ"s��J	���]c"Yy�b�/X������Բ��˽�1���G�BP��A9���f���Y˚3�A��y���E��mpc@r�� !a���v�t=��A q��ۢv�_a�P��=*l��I9 ;����k��@x�����=u�{���߭BP�Lq����R� ~�3ƚ�%�0O���jl0�%V�~�i�X��Q��7:=���c�?�89W�[�y��O��U�plV��5�#-��4Ԗ�Q�h-n[�jK��CG���XC���d��Թ�  ��IN�h��P�$9��^�&m��Y	�D��i� �lBxN2L�a���Dtk7��`su,$�=4UāDlm�6�� �)L�^Ta:��M��04-��>�҄%ϴ� �w��B)�;_�jD�*R�L��!!϶�gFr��1�f]H���~<h/�i.��@���~=���L,�=�Ǧ�� �b<����H!�0�{�M�2*�5��X,AЍ�����-1�w����|E]���	cF f?�ڴ�
�L@��!�)!���<� �D��1����!&B��,�4IL�f]�O} �� �H����"�"�^����$�J���3:
^Ȫ�� &�mc�RmN)�+��\����FW��t�ޕ1a�~��{�kL.�oF�6$үX�Y(Q���
ē�y$nR�&n<��]�ڒ�1_;h�IS�յ�s�� XI���V�*P^�1�өZ��$[��a�P��)o fb�#�����I+-A0.�[��Y�[q�P�r�h,ܲ��l��#6�Q��P)l�QG�q�0�g1xs�b��8�X��Θh�C&Y�{e����A��zҢ`v_,��C�m��a�K�E��̀���s�@�b"^j�m��T1�����0��NO��Sr�_�t�� W}��w���&���~��4u��#�1t*4GBT]�(������3�芉���@�=�i�8���%����� 5����F|�v
K"]����HJ�ܙ0�� ��&�en>壍M��'���QQlB#(�-���$���w��:�#i�?ɓ}L�P��2TٛΔ�C$X�3�y��4�3�r�q�� �2=^��P��ۇl��Z�1���:F�D����Qd��{zq��.'����,L�C���3�m�0&�y��q;IC��B�4��JCH��6�]�:$Yp���CC1+�>���hT+$e�#E'�I�S1N+m0�	a0PDK\�H���!n�4�heu��G����p*�2����<))7+m�F3;c1�Pdpb"L��2����%\��ͺ#�fl�m�S.4�
��`�O��N�M9`J��'x���52�e�U>vnt�mC"n"a9�LvU�ez�4$��	�z�0�n���S�+U������x����"W8�th :Ǐ�t������1!3o��@[7��O���f
%;\�z{�@�+����P��<�σ�:Q ����ZW��[��d�U�TPZ�/�Ϟ�U� UΫ���?f8��I+
1lm�c�Ѹ$���M�fH��m,&S�#�
���ח�H�*Nx����@ L?�mfq�T#n���&1���BRq�F������5�4 ��	e���� �H9ܙ�w�έ!F���1�D� ������B���I'��2Wb;�jXH��u�Þ��V�Ly&Y��rԜ��0�`���,������!g�:b"]���WM: ,��"�D��`a���dpeD��D��H����'US���ղ[4�� �$Y8�+3��D�[SU�/0,KW����C�T�h 9ief�!RK�
�J�OR��)���$H��and#�!���J�i;��WB��E�@�"ڪ�H*��N/#����T��R���
4�$��Ä�m�вQ��iHÄf�����d����^J�S 36��0S2$R�g�oP4��w��<?����k͗�sO1?\��h���y͟���
&���-�j���OT��/<N��&�Hc�p��BTg�_0��i"��Z����FD6#	ΐ!fӼ���$qf���v5���f�Fڱq��	�Ob��h$.�cs��=4u(�If��=��d �JRJt���Bҥ��k� )�O;m���Ms�sn�����K~�W�2� �g��=o[��g1�mLe��&�W8��
�p���,x�%��[��C�ZZF^D
���h �ߴ�� ��R��`��.���S j<�(��צ4�(��q�GI� �����2�MO�?SӯM�̙q��h�Up/���ґ�Ȋ"�]�8҈HU�z0������Lћ�j��`K`�c*��AUfg'�Ye(�ܽj�������H"�$��|��D�KbX��Hۤh��V�jMq!R®y���5�(Y/g�gJ
}*�x�g,�H��y��J uu�)�mP�o�� �{==��Q����:��ap�1���oqD$T���*�Bs��"3SQ�X����#tV�����"��fqF�
O �+�Vne�F45QбF����N�)��w��)�a)��3���������G]�D2�;s��;��6n�	���5/p7������n��X�}u�FN�x�s��Pb#؈�s="���d�&HN�/u �ƈ@�_�άL�rE�1%��Ҡ0���E�	�r]�+��n1����O^�ZP����1�ƈIb��b�΢4��-�g$ԅ��X9�oB3N� ��#5�(H�حڪ,ZU":��gT�,){��v�F�M�BD,Ĥ���{�0��y��mN��l%�%L@�i	�,��oh	 H�"��o���VRbK��j�:�@����I��牙���j}$�ڦ�:R�:��Cx��~���2xܢ��RLF @�8<+4��IÄ�)�/��$�nbR��$cK\&��7��La�t�PYL�ؽ����L�bg��fa��K0	�$C2���� D��{j6<�7d��&��s��$�FQFj�TW���#id��������i� gL�2�y=�Ȁ		*
�H�s#�F�,�8��d "Lm��!)P�L�.9����X*�7gm=Ed��(��=΍�U�e�8�x侮  �S�~]%9��$�����9%�;.&�;$����غ�ƀ��fҙ�|"+vt<'�FH&� ���u�6o�J�,���w�\hѭ��fH��S"u?{�� Ҁv�C��m{�9`�}~���J�-��>�k�L�0�Ϙ��K��,��moUXH4�FKsaמbt	I�������ꥑ;'�0��Z0�����ȳ�`Q�,��o�Ou�8�d޶���Ұ, ux��Pİ��(X|j�i�-���T�%�X_$&��ǆ]�%\�gK�aq�����	g��t�Dϣ��FM	F��]
 K��B�Μ�K��s�Nם$�e2�}�Ζ��%'��F��cw=/fw��X��pvg��� ��7��.��Ճ��%)��i�Dm��n�F�#y�y�}@Y�cn���M�Y'&��11h"!������NY>Vt��Z�0���|�hsq;c�:��%Rm�O|�)(��f�_�u  ͭ�ۏJSh�"YI
n�K���E ,R�~�7���+|����� .YV1�gG���:N�pU�f,��C�t�r3����0��V1"`��k�h`a̰��&�9�� ���6��b �41�!���xv�	��`I��&��� h@i�ߌ�w��A�q�7�߶�mRM_|�"B�ȿ�m_,�K,��������@ͭ�m8���X	hd��\��]H��4G�bŖy�j-b��ДP	�b$�C�N�YT�r�q�#~-3"��KЂ���Ǩ�ӀdLK9��~󩈄�-���ԇS@rn�iƆE�Y��s�Ϧ���H���t�Z2J��un9��5.�"�3'��D����ۦ&�� #�R�����Y$������ӥ��L�`d2���HA�b*����cK��R䳜ę�Qc�A8��6��hPX�.s�z�<�M-GmŨ�����D	�4��qI�����}��-��m��.��&��Zԉ�3/^9�oQ�K<����o:��$I����8�bS��#A�/�X���U	��9�]*6IM�����g��b���!�I6�ߞ���X@�qȗ�@�Fry�$L~tP��z��!
�2����ST2޼s��#+��h��^��as�����[�
�l�{7Υ�C�(��}��b�u!�?�R!e����ԉ�s7��s��e��s��Ι*������J�g�y��'�PEVm9����	I��Ò�u�W�����NB�r��?֔7+J*����:0���[�n��X�3�q��t
 8/�ƥ����46f��D?|F�$�S6mƅ�w��h�fuڟV�=�7����h1�����:@%+/9۬V�#)���d�f;~yЈS�y��Ƅ�b߷��}�$��g=b��0�Gz�P�濫$��j*jz&yҪ������"	��Li�K	����������Ǚƚ��*��nw��ҙW|���Df�ۙ덳�ñ��J�� �FEM*�_:s

�3�����1�Ne�x�&�8��8����u�����Y� �w����Ag��g��E &+Vϛ�8�*�6����@�
���=u�9Ԯ�q���a+8�䨺��7Ǿ�}:i]⢫G,���lm�@%fX����v��+����)"{L{���Jq��Ǎ.@�m޶�g:O&g�����v�< '�w�:[+�L�3����p��=>�t ��}���Ӕ����B��|����e��n�W0Gs����s�1!�Ρ��=e�����L7i���u]u��?w��=� � ==��x��	z���u���q�!Py}�~��c����2��^���}HM��#Θ�1��:� "����Iǝ=��~�4�������ΐmɺ��v�?��߽� ��n�/��	ʳ;Kbd��i�`�lr�o� ���o<�^�1Ω�C-ʿ�� �m)c>_�8��Z��m޹� w� �B��^�}&Ik>=�L� ˄(T�'߷�As��1OmIR�.�� Z���O��rdo����Ƈ��ƕ���V[]$	���0&�������I��&�������Њ�ci�۩���;��������t
!Y�gw�G��G��t�#;��[���u�:s�����Foӯ���/~��/G��'�1����0H�ff����d�"2N"6�G,� {W��
�m����Y1%9���/�Sv�����2��b��6�Q,)�<�II�I�#s�p��Č�61��Ȅ؀��q�y2�[S�<~|�lV}��ﾘ�Tmq���H�zze�ycI3 ����ގP%���hg������.�hp0͐G3�f�2=o~#�e�K�R..x�q�+����!��[tf��` ���fө�_���M�$��պbD�.��K��%Ȝ�5���$beƔj=8tP�OH��x���x�ڼif�'=��w|g���85��޹뤦F$"(�@�F X���ԡ'e��&띴���4����K*P��sD�t~��	����Έb����-�j��$����/�;��A���v��n��nc�ޢ53�b$C���4:<͕Bkԃ�\FXL��ǥ� ����O���� ůDN�t�*Dر#4ɒY)%%��"��Vt�!&�I� 	e��ZP�ő��[�~BPD�Zi��I��6e@&� '��pк,������SΈ�0@��B�%�c,�D��U�LN3�C�(9Xb1f�i[Cj��;��D�}>���f(Ǥ��~�EI�c=*������-tBQ>����y�;m�_��%ؘ��c΀�Vjag��g�.��D �?�m�e�%�SJ�=���%���M&n��z��ٝOJ*D���H��X�5�&T.S;UV��dܑI�=+U�*,8���޳!�}R#�񤺉{[�ns��a������i2�b=j�ם%I�v��g��߰H � �Kw���ɂ�N��z�?���oΡ,��&6�<j�$P� #�A�H �P0%  ���T��BX���V�FZN�� H��I�pRE��e
�Y�/��4�eZѓ5&�𤝘d%	:3Uu��9�PƧF�Ѕ��d���t־$��h�'Fӌ�%$=j���)U(\��Q%�C,�Yފ����������)ʾ}���&���l���NAt1ۘ�E�:���qy8�oF�Va3�o?���B�rc�w�OM
A������y�UhJ�-���G.��0�2��b�KGnE�/�LV�2������X3P�"	�	j6�H��6d���(�2]��m4%�&�}�(����7�]]ai,�"~\6F����}�Ɛ%Y�Y�k=?�`����t��'D�4|!�B�K�yΠ� K(���@�8��R��X��+���D�e�]��	��(���&&��a�j|#�d��h��FKX(��*b�,��N� �nƑ�s�Q�+yj$�=Ѽ���ƦA �� ��o��|Q��T�3 ��ዜ�f=:��� � s�0&G����@D�w�>w���^c��3�� E�1R{�`�l�\��gFeC� I�q�R�8Җ%	?q�6�t*�g3�_�Rg����d�"}oy���eb%LŦW��5��K�>�a!It����)� 6�!E3;�Ɵֲ�I���K��T
�r8��o���1�V��G0�!	����2�THҐ�}:q��)�!g�v�Q\$�mb	���NJۺGN����A��Q������H��Q��c�?{i� 8Sa�C������Q��*"��J�CR�b�%�$.�A�:XD Q`XV�1�ZQ����(b�QbA$.��a!E�y�gX!
��1�WWS1ac�'C��T�r�wȀ� ZVԉ�":8e
��G�I%�ɕ%AܒaOA+�	%tr���� �"�P&t�R�$�E�s{Țҭ��G��Rc���^��_wF��P0�4U�=ޞ���x�� ��F�Fg��	ޝ�	�sǌ��I���I��wƦ�d|}<tҭ]f{zRJ���o�ƀ������oJN@�t�38�"�����;�z���@'4�m �_C�:ޢ
ٔ�޳�6;��H_֔�GU��eg�M B{����/B����?����<��L����΄�_�r?uS�8=�zL|h��۞��`�� ʆP�h��Dʦ��{�<�Ed흊���̀DM�
�b��`����\��R�D9.�MI�9+���G�E �X���(z%$R������8��]���v��*)���Q�{h�
�U�4p��7�����T��E��^91@YO,�h�a�z�`�Y�x���"FH �i�ƙQV���g;�^��h��2�\Wm�v4`�� _�,�'��d�*#�;.� �,Sq�}q�;�sW=��[�lq�m(gD�d��d�B.����D��-�?�RT�DÁ�����cJ�[����i���F�6eϒd�+�g�+���bcJgsy�TgP��\��4�7�T܆�	��].c�;�;��ܬ�3���o���3ku��;~��(f�����Fe_,x��5�tC�����lgN�����Lތ:��nW�B��q�X�2K� �},ݧˈ�Oo]���)�|�ΪC�O�e�?:`Ȉ� &�b��W1�����)�k���HY��ۮ�09�����*(l�iF6��)JW�p}��ߵ�^� �
�/c}�����W~�A
f/��3�������]�rA�k���H��cq��X�4�	����O�j�#	��L
�v���lv�|��̇���뤣*���jRPLr�徻�SN����P�]M�E≾9�}���$�7�>�����p���`$�&߹�I�����n��)$�!'��^������Hz��bzhݗ1��ѩB1IJ�;�1e]���#���Bp�S�v�J��o���	B4�|<���q�j��s�݈�Du�c�{j8[b+�Ƹ��;�W��΍�w�I�"�	m�:^�
z���z�mq���^��F����/����Y��v4\6q�1.�������ހ`)�_ם[��S���I09���u�T����lz�>���@ۏǾ�����t��S���WƕNC5���:xX+/�O~�ixI�%���m�
��{O�F��lif�c���z��W����|w�g��f���((;<����&3`&9��<�В)���M��3���b��x�8щ�dV��;�"q���J�S;�0^��
ɜ�A7�ր)��{�~��"	�4����<j�Oޓ��s��:|(���a���ZL̍�N?�h!eW�Z�Բ成�����q�[VH���˼�`8�w�ö�W��� {8~�u�J�!m��� |gQ/�]Z����_�����HH�i3�N�v�_ ���7���o�����@R���1���������z��_�϶��}�� ��zxs��������9�b:���SbD������P�w�y���r��~��"�
��~�B���~���ί�Ρ��������������t��/�����ϹԼC�����������^=���~4��'jƁ�-��c��u]�f*���� ��L�o��gE�&:0ݬ�zV���&b����0��������u!3��3�ؕ��7�2i�P����#�7���<ic:b��f ��߶�0���I[nw��:�oX�@P"$���7Z1�$e�fz_5�Ԑ!E�^�^�� ���3<�"#A}�Lر��ߗXpP*g�n{N�J���䆤硳�����_.���y��0r� s�� h.{B�m��2i/���y�K[Kޢs�3��m>��*u��:�I���y���4)�f���
�:}��oΖb�q�LF6��o˟�;��2��EX�߿������o�w2�h�o力��v�.6�1>�v��W�~��������Z�|�����Ư��X�C��������������Ƥǫ�������gh��i�S�!�P���x�9��94���Y_��4�X*�b�����=��B22�$�g�.@u���8���`��|m�:ّ+E�|�j�W��ATLl%d��x w~�?z�Q����L@3R�����vxbD狆ޢ�Hz�6�l��U\5SK_��FB&y����I���qO;m.�b���N�8ŕqMF1�(Si1�Ж)��š�ڷ�T�2��@@Ic'M��EX�����t�'&��$�
cO���I&!&�&� ���tp*Xz��*]��'<��֝�E4�ٗy�{R�U}���
T�c�g�hq-�ػԼCk��ө3���󠶞���=��C�5��&-{�}o �=���Ms�k�7����}��e��j��I��>���gPly���
[��D�=��<��'����|���,<U�!��׏�� �Q�� Ğ~w��ڈ�I��=��� �;}��Z)��m5�=Sc4�
c���e`Ř?<u��E#Ơ~��g���u�׷�ra� #C���35��� ��tԛ/f���a1�U��ʡ<1yoB�����jY'����@+7��ei�3cu3��i#h+V�3��6(�2Ġ����)�W�!��l�Ӈ1`L*[��gX�ePH���7�1��� �r�m���T�
J�j��|IH�scLK�H�/;c�bi%��,D��M��!0�=�2^���!I�\�g��0�jQ���~�tS�c���t!"���M�k��>�5/��ԙ�W�;����?�z�Ӑ��
����ڟ5��0�Լr����ܫ����� �m	x*�o'�T۝ݣQ�_�vԼ��SbU�����@m/��M���]����$H9���5|���_p���M ϧ�� L1^�x�>���������w��a!	������� ���\�W�`ל~k�4Ęd���*ޓ���܊̻��_Ƌ8�&����8�?��9��:y!��Rf')f|�#��\ZT_����R(�k�0���/И I0b"'���R�!�'$TF-.fdL�R:���P�;	$�~V.gI�&%��曶������͑=j4���%J*Y�p3��d`���w��}ZEc������)��� ����s0�s%�9y�w�pi���!��\ND4,�h�^�Dq��B����^cH���5X4��pfT�(�1�vH&+VL���*G|���:�
�,!&�4�(��=;m��Bǀ���w��fjP��ҚI
<.��KYC }���IH c13�z�q�A��'��B/5�X���sl�(��ʻ�CAT�ə����v����x���lJ R�\�Ox�@Ƭ��su�	��V�s9�wh���y�"]�X�w���TJ��!{��q�II�6��LD��Ү� �o��F�<1�a3#�^~t�;�~c�54��c�:�:4hL1C��;�:��w�y����Fo�O]m �툣|��M�XrN��qeP�"�!:t�Z���˖{t��M6���}��������@̮dM0��NL��hI|�+9g����Df?|ĩ̮ۛ\Tw�Q�L��'m�Th��^��h\�I�bҖC����@Hd������ A/,-<ٙ�}'	�'�L��7�Dd��j�ܱp/4��F�3S[���j1Ж�.y��T��|��{Z��Ζ!�D�-(j`gH�X!��2��+�D�i�ߝ�ЂQ��R^�,%����J�7.gV2*bX6:s�g�P�aF\d^��!AJ3 	 �$���5{��=�1�z
��h��� &&	3+WN��6I�{
L�F�\Ćf�9Фe�M2�:�T��f!ɸ	�⥖"P��}9HM��ҭ�vW1^ɐ(�/��҆�`�J�x�-ɀ�ޱd�پɄy%�C�� D�fU{�Q��$������:n+�e"��v�-6�	��fMz�x�F�EvK�F`����y$��0A<w��@&��z�����1�勞�F�K�;I�@�оu�����+=�~�O�.��}+�Q,E��բ�t�0�o��d>>�j�����	� �o[s���f�6#�s��j����=�"b#�3���,}��E��*��;lr�h�\�g�V�����|v�b9��Mz��~u -^� �3�-�E�x��:4��(P
o��t�X70��u��C򴸁M���HЀ���^��ѪKD
�c�x�p��X�E��񣒎��"�/��j63��1�#��6a�&9=���+EU��#������+z��4l�rhZ�7��f"%�yh�
�N�i�Ih�`�(��@$�T����KA[���`��")(�"��#[*z3s;(s&&
pK)�&eY���0�; F$�Wx}�f%��5II7�V��d��g2g-�:�(F@#v6�bԌĈ\ak�:)bd�lX�1����P!mc���gM&���CNn�E�
&q7;ri�DJ�O�CO���XSe=b7t�
8dFan�(�LN�2T��ٻ'w��	
 ��|��А��y���GQd%4�ǧ]E�(L��Q�ɁG`��w���Hi��&p��_SHF���V�U�Mg�_�~��$YS�d��]q8��ȡ��^n�'��*8�c�_�?�˛�F��Ͻjem��Ͷ�K��Zo'U��\Υ ������,F���֑9_���I"rh<o;툓l~}��|��i�F�����c<�Yt`N!�=|�Hu`��]�� Uܹ/��w��E �Um{�/2`�wYl��Ӡ1:�fg:	�Ba�C��� �ȶ�f7�F�)H�}=��yW)��\�Nj<�r=J�s#Q�:^$	�&{�D=�Bh�)X���s@LD�ó�
N�3��b�,�����)a�a�
S
8�ƔƄ�yE��ˤ}ȪF g�ةuT@(��1]r��-�X���Y5�-E��f����)"�%!�^��"� � �w�W	�M��f�~%�!� 
_2���"����Fvw�i�eo[U�:��(̌D��4����M����L��,̸eq��jP�8���O�0P1�r;�h��4 <=c$:2M�6[H��u,I��܎�u���ČN�1��������Üޖ��\�3�^��D�k��u�WRgш��ԡ0����K��x�2�/�l���:#M����i���(��0���a�N! �� c����'�;�sZt�;�M�i��������)s2�o5���Y�� �����H��?� �v?7^6�{��ve�WX�lg����x�Q��>b��!(Z#��4��i[�\}�P��|�	���}N����C4� L@��28�sP�K�#@_ Vی�34�c

aR +88�ӊ��ݱ��q�9G(��H1�G���R�)�+ʬ%�����r҆�nz�Q@P� �{p�3i6Z���:�ĸ%M����Ԃ(�d�,�|hu� N�Y��t�$&XKq�Xx9�j�YD��)f� ͬ`�����T`��Q�&.b)�͌���'@[.B����ӹ����;V޼�I�����U��������s�oLUoR�"K���G�� ҈���ǓKuRžmN�t���Y��m٭3�2����P���JǼ�a�q7?<i.���jV".� �� X�D��[���v���S��8!�a��:$���;K��o�!,BORJ���H!��k�5YD��ӥ��
��q�O��d+|�t�@ÿ�M(�����g��㾲q'���]�k�o��}u�+�?�d =���4������Ky��4������D�q���u��`��)9ɍ�Ί�U8\u�Ѓ��%8�dNM3���(-y��x�&x��ϝ"�7��`pD4X�R��%�����ҁ��e7������M�=fK��-�r���rg&�LDڹ3Ь�%�`l)��\�3�7ʉ��t���6��[T衑�W1�����5���/:D�#b���bD9vم��D��W�Y�o��A��H�|��|����~��ƘA�a(�|�]ט��խ#��:u��˩1��>u,v��n���~����z}�n�0��P
Pw���>%���I�ē%S:��C*�z���_��C*��f�r�4)P��w�}�-W�%s<{i˷N?�W�� ~4̋���4���+*�Ӯ?�l�����^4�%1�� �����Go�s�հ��u(}���wU���@A}[���֩r��3�Wz���2���V
Ŋ@�-��� !ʠc�Ît����p����O
(curj豺 �ai�5���̴�����	 7QgPu0��V�&�'}U�hk�� �F5�NM�s:��?	�-L���#��s������·-�@�L�,�Ǟ�#5��WH�VH��J���� @�MOm�|�韮��}�� ��=:��h�o�P�~}4L�����������Q�_��� �	o=�Ʀ���� up���Bś��ά8>ٯ����3{�qجq�' V<�5���Y�)��w��	c�>ތ�i�g�k��@� �l�o�t�u)�q���}�[�i8����~P��ϟ�f�'~:�j�j�-�l>��9�~�� +e��x`�o��A�����]N>�ti�lk�v��He;o�����cxc���_�����]ky��IJ��$�Ds&�gI �`*g+<�z�@X2Bț�c6b/S�l.J�-^�B�eFy��mwEj��K?h6v��	�9��gEb��[�8�����D��E$�a��&�����#��v$erm�p�4�6e���B���$\"f$P&@H�"�i?pA��=t%�椋�{6�L��&$�3�
A�(J�,�$��]F�ZP�~}4����}�/w��Ԝ���񠶞� cJԒ"�i?��9p~q�o�W��p~ơ�E��~�F2��/��Z'@T���zFeC��o��IHL�?&�4���O�� ��^o����L�����d�\�&vgB:�����#	*M�����BdQ`h�	�NƓ��\���WmM� L��]�������̝��} ;}�� ��-)�v=S~�������C�X���Խ����닖NU�}�M@1�n��U��������0\g�q��m�G���i�6���Ƥ%P[�{i����N~���P@l�O��X�����m���MK�r��������o�]�10/2����50�nb���o�Dmӥ:�Z,�,���BSm����B�'pT﷜�tq����;�I����~�D�7�j����k!��P#@RT�|Y���V�=_��A��O��P�&`��u�҆]/&޺������N/A��!����U)��A����M�1;v�X�A�qaժ�4MHP�l�]+�427ox����L sZ7�:����v����"�/1?';��L\}���HZ�<F�?��Ɖų��O�#BR��J����U��`0��P0N�
_}�0uю��W��LY�]�za�@��\sX�z�k;}u�Ԩ�+���æJ���i�UYX�r�㩩s�C�y�M��Xw���ceqBS`�`�(��N��_�5?�M��\�s�r�g/\��BG�]MK�VK���dL�g��R�M��=6��h7��ރ3,����Q	vD���xt��[�p�=���h��¿}{(�G�o�LE���_O�u",M��+Aa��
�{+���,C����'�T���d�5� ��X�(��VB�<��U�+�"e����WB��ITK��;N��oA���9�����:˹fcٺ��#�"g{)�n|N#��]����X�U�rIqe���v#q:s.� �
 �����Sg$�a-D1�5�@�A@P�[�{@\���Zd�a$��פ�j 1/ad�"]ObLA�Q2�y�1�4IY�ʳ�̆6�)�5�ydh��Mvajz�5q�?�o ;�}kH���KT��� D�d�����q��yA5'������N>��He]�	�n�nZ�]&��!�5p�67efq[�V��g��Z����iDf��Ǭ�����񚘙`|oƬ%�g��z��ԋ@�L��o��5�A,�B#2^�Sq h��X�G�:)AL@@��ՆC@9"��6%&٠8��Lİ.�=���=>���@�~�h��y�/t'��OY���J�;�&?:�>�=4	��ߍa����c��	㕸�g��H�my�c�>u?���A8|uӢa.fMö3�C)�'2�NgK�%`��lB7&��3bڛ|� ɰ(�B�pHTUY)2Ub�T u���n� ʛVcm*fh6�t����߯���;�{�6�m-f6<w��
��a��J��{�y��K);�n�=�P؈M��J��  8D����&��A'�5�bF��� FY%��A���`XY����@>� ʐ@�.cI$��Fؔd�j9��j��A�$�S��x��V��bM��u`Y���|Vt �����>��x\��:�1��#�>���	�
̟z�1!Տ�h�z�����}}�0G�BA��77?���]�q߷��`Kg|��A��*�ϰ�����#����Y.YY� �*&hj�9h�p�$M�n:��>���W)z�8��N�H	4mA<aK	���Q\�zv�]��w���ޠ0�2ƒ��J�C���ӍPt�m���!�����+�y�X7y�'h�+Ւ��������7�~�^���X�E��McR�u �LA��s�1�e�V*aB� �(���I�]'�4iH���c����=:��k1~��<3�(�}
�}�b&�=1�R�z5��%	F'� V~#�mv{Qw��]H	(����tM$YkA)�rh�xHc�M�^��F@!&����H2����5ZEehFI&�S��$�eݘ�U4+DVX�
�^t)��ѳ+r�Ox6D��Zc5:q)bYΌ�x��翧Φ�q -�w�J�d���oj����7X���9�Nˑ���J�D�m����� 45��˩��7������{� �i��j��/��.ي�[�{je2�=6�?LX�ǟ]���c�����)[|�M��DC���6�W�΋�a@ �&l�Q�h�2�lJW�����ܐ/p֢Cz&e�e�܍,�%�u���Rc��|�X�����/߻��#O}n�_��mM����N*t����9ƃ��U��c3ZP#�=\�H2U�MF��#k�w��2H���h
-�� �+�c���))��MLG��S`%��J� F��X���q:IM �^��iQ�9���5`��s�!�h��GJ�DC�o�=�G�?s��?zN���ί���:`*�S�L�g�6� [R��`��8h #�qn�}s'���۰�@�iG02pp�;0���7����2 @J��.�ғ�E��m��&)0�b"&J���j��Ѳ�YArwG�&��D���n.�o��8>���_��Ru:���s��� 
�/��xb���_~��֦2��q���b�}��ӚIJ�'>l�P����7(l\�\��gž��P�X��~gƘ���>����D�����%���Ǧ�d����xөb�c���EI���n���L��b&.�ђ�kW�Q��oe���`�H��8>5,0ofc�ƫ�[�f�Kb������~���:i�/Sp��~�5p��OΉf~���A@}�:��kۧ^��*�{�ނ@���̤H����خ�*[>���� A$� �!��/O�A@��.��$ѹ%�؞���mB�egsf�EV��Q��ܞ��S�L��?�^MI"ߣ��Zg3�̼����,B�O��ޥl.{E�47*���j&���� �j;������<t:m��fY-'����4tm5�˒ !�*��Ob$�CbBbI��7��sNc'��.F�Re�S~�5�6�!;8�#5<h!�����{�H�`�E!IQ1ҵ��SN��ʈ��ff�F�;4��TVT�1�.Ħa$������"Yl�36��9�W !�+�槍M��Q����c})�y�3;0d�_���\a���	��W��JT����Ҭ� Pmu��J��eU4x��SbS3Q�}|�t1k���ީ��X��i(m�6/� !�_���>�@MG-Y�vvh�ܾ1���=�&�4GJ�w�q�bW�����5�(_C7� $�����3|�=gQ� d����7h�_'>��Gns==zh���uӖ@>���D���������嘘���R%������b 5$�
%����~]�z��jt��z� ZV 6���}� ��3w�B�[��j6�E��~�����@�}�ԂD� C,,�Tj��3�g�:G\���iDD#5��Y3�㺯�z� ��y�yǎ}tv�ěܗ8���BD�f*b}�MG!`��1�~�Ȝ�+6�k� �!�u7I�:1&B�2��$Τ��
�@���Ȉ���+���+��5��@��>�5������������A����m������ c�bZ�ƒ��^�O���u'+�}�h.�5�4�.��+��  ���}��{[��<���1��*gǮ5�S�e�"(��Z	б : ����
6�'�Q��@��:U��k��0��"��
aLa����@��Ϧ�$D�m�gI؟��ڗ����i�IaL�3�\�ݟ�秊me�� ��s��}4X��#�����m<�m�P�%~� ����	sߤmCq��KE�6osB�.�ʖ�"��`n(�-_:5+V�38t���K���~6�'�JUo?6�zr�u� ~�L���m�ݎ���9����l��y�������-�.��<G�RcIu� r���ԟ���P�ĴM������fK���?ְ&v��Kֺ����9�=I�>��B�&�\y���K�N�tn�ޯ��_�>MR��"O�U$gA�TN
���К!O����"$;��V��H$n���z�h�q8���C�}=�@E�����	O/�h���7�f���gƜ�=����E�I��{�Γ߾��h����Ʉ'T�����������ev���w�}��3�Iɶ���C���Ύ�/洲�gu��v�w��m,'���|kr� 3|��Z��R���U v���?��f�0q�/wB2D��w��N$�ě^/���"ı�c���J��F)�������TY��y%�o��}D�Tt��
��yq.��`A�mv�����D�n71�:�lpX�"�[�Q�xG&�J�OY+Rl$h��yϝ"�y"�p�]Ng��Y#���K�t*t����mH�1�3y��ֆH:�㓷Χ��=��x��DF��E�� �(����g��1xs�Z��e�=K�_I�[#�[$ۗ��Mi3Xۅ<���Z�.6��&��BIܴ�v���!$֌����H�,ɨ8s�B&�����/��������I������Mmu����<L�im ���"f�u~�Ϝv��0����Έ���uҵ�x�gYfv3���4�\zէ��Z��i��f���]��|��	�/?�u�m���0��`C��HO��\q��b{��
�Lw����-��s�����t��j�����.v�[�Υ�	1�0N���ҵ�<�y��u.}��Vژ	���=��Fp�87?�̨��A�� �=u)e���*w��5����`Ʊ̳'Y��o��Φļ���V���J�b�h����(Pa����ɑ�qL$l������V��W�M�/�: C2�ǘ�.q�FU��{�$x�$@XŝH&�*���a�϶k$���cfcy�+hp871�����VK�>jʹ��`�RQ��;^��%�$�w�x�F��(�5��Cf���7�H�X�p�HG	N|m�ѐ��l����տ�7q��#��r
PDԓ&'�h�@��M�ǤhR@�$��H�&�GF��A�����t�iC�A���z� K�0��z:@��`@$��6�gDZP�� �#2ytĆT�Z2Í�4zgbC@e+�6�0�	j2��̃�U`ȭ�'�_k��l!� �bwN  ����h��Jd9��qd�I����B�SC5�n�ґIYNŕ��zPG0�����I�r|�ʨ��N%��%y��r�)M�`^�w{3�[)0�(��>�΀*�FLX1Ss�]HD���K��?�f����i�B2�G�UF*�f�b�d��Ƌ*S�8��ԲKp�	��R�
WyE���V��;c8�z��uyIJ<������nE*r��̛̦��.�5-�5~�ژ\0�!�����0�1..w��"�.�����M ���|�cz�,�D��s��cmD�l.��nziG'�4���}1��T@�o+�r�"-���ȨK��9��}���fM����ϊюQ-���}��pf%�7;��1�QS(2����](��0=3��$$�8�0�j@��19�i��J@	���Ż`�@���6x�N���L�*��	�8�M�~ڀP=" �(���8{V��Ve�q���W��ψ�=~4��RTi���|h� �`l��l�H�0H,�1Y�5
2e���o��E�759��� �
z[agy�SRe�<���w� -�@R�M��md�=�lf������΂R�a.���f�����*�$Cfd;��u��;��=�c����AYe�os:v�$�7ݶ�[1Cň�zh��`0 ��39\�f*m�sa�C���j#����;``day?ez�f�s�V8J����K-�85'�6��<^�� �	����u&�dI���uDr�g�a$V�K�q~�Nm��,D�1;ef!3�{iv��yd�"�q�gTu*��m��4�������n�	����c϶5 �I���G|gW��
;��j ��Ω�{�|][0U;3�b��"��[�0�`);1�4"F	���3u'Q��eEE�G]%���Gm�LH��~��cC�;g�q�g2���Zt$^�\�7����MP��b�ä�j7=zy��I{�5/w��q��I{`_�F��{��������BA��^���� ���Q�V����cz�Js��!�&���B�S<�
C�uݟ}��h���������_~�� �@|���wK���ߎ���,0V�{F;cQ�-��u�������g�&N�)f3'R/��qHh"[�u�S���N��@&
S�c�^���LI�c���i�A������љ\���18&� D0v���z���ϯMFD�Em�}�%QDҎ�Xb��������\V�����	�?:FV� 11[�ݚ�Bv���T��sИ��̅V��� ��Jd���7��C�a�m��� uˌ�����D�����DP��]��,�D�|���F����b�9xf85�f���+T��&�A'K�Tf}cMA!GDn��P �@c�F��y���m�F�@�jӆ׷��7m�� ];ޠ\�^�=d������l����0!���4�hE7� ?�PŢ��x@���7q7�38 �A��w���8ǝ���1�mD|j+go��Vw?Rh�	���I�[{m��e6��GtdX,a����1�Lel�����]&~Ѿ��4msQh���3� ��7F�.2��i}=���^1�p����a���ﶲw>�����F6���y�>���G�{m�����q0y�'�m3���7�܋�^ci�k�M���}��@���O�C9B8��4�ݭo�||:�^c��ڈ�\�O?f9����g�L}^5*Bf�^���1�5$�����޳�͌���;F��I��Ϯ�8�o�mv��ĵ�g�m�Ό���xԲV�U���g@�s�N=9ѡ��و���;���g��3��Q�\�r�߯��MBB 2�dS��#�������ƙ�PS��]9��\�p�_�o���z~�C�v� u����a��1ϛ�q�ϯ�M���� �H	dc���~�	�8�%}�6�y!�&oǥ�r
��UoF��U�޾�����S�x�M-���צ�dIᓣכ;須/������)��v���7&���}�f�'W��Ѝ��r�﫥 K���v�\�I�X��e;gD�)18f}�Ε���p�u�x��z�o�%zV��0�Z��6�G���Ǟ��@������}�8�ǟm���Ƥ���}��Cu��Α�f�Vo_qQ�,\,_����1�����	�Gfk��v�R�b&����(�ާk����mF�����m���
^T�"����zS�EL}�oT&9}������ U���Y��)�s���gD׍���?Z�.9e��:n��*s`�=Y�6iZS��K�N��9���/A�B.���#Y���0���o��y'DC&s_���3/j���Ao�]
���(P�1߉�W$,.ѿ�:Z��� ��d]Iޜɣ(�#|o���*Fd��U.�1��VX%��]�Ra"BM�� �ɡp\��T���ƄP�z��/ǝ!�� �3�uc��߻i�P���{=>kc &v�#)ӷ�]
��_y�f;�L=��2r�O5��F��,�v���=i�Iq���ήwm�;��;\C>��Ι�3/���f��V�?�^�zf�3W��}���� ��}=��?~��2~=q�ڶ�JX�E�����Vy�X� xtT9�����nF^�&�����~���i7��t��C0�n61�x��M���,�=u(M0L󾟼�W�{���4ڰ�ښ�?3�>sY��o}5�o���hG���Б��ķ�ŧ����Q�B�v��'A[���������i��J�C�����^6��B	H���t\�����rNz�B1���!B?d1��5�9?_��� ~��n/n���JH6�w��� ��H��߰�a��+$m���d� ��1Ơ�m��Ή8Bm��;R�h��a)!�	���L���DFn�突�������x�@(���Ѿ��?�š�;����ZbbC��BG��LBY���n�;�Lw�홍J�1�AN@�
��Ƅ�� D$)٭:�$����(��/�=�|�}�f,�,��������b,'���L	ޫ���N��$��s���<c�&/�㻿��u��O��Ὢ!|gOO����T��ϯ�ly�X�խן��]3�y��� 3����_�4V�x� �_=��W��7�q�z�΀YK&���e������4��2��4�}(�ﵼuC:d���Qܡ����Qh0����y�y�x�J\�<�"P�Q*��<Mj@��ҺW���U�������_Iz� g3׏O�C9
9��Όa��^�|� ��y����a��{z�
R��1�N+�(B�K� k���H�"6�!�t��⯞6���9 �<Z��Κ*�>	�2du�fXgY߭I��y��>�� �2��t7��*!���w�<�A"*y���DN��Do��D�f`IT�I^�h����B~��E��	
A'^7�,G�w��=��ZL�u�����p��<��[GD�&aOM%HX��}魩����: ^����E����l����s��|iǒF"��M��O�0�� �5����#O��6���;O��}�`잽��Tg:�:�q��N��a��s���������$|D�q�=������R�&������n�����f���?;N�����3���.o5�]�프�B��q��:�@=M��s��'fDX*�;��t˚���j�[e>q��·if�q3��T9Ц�[Yyt�K���ey$c�ߋ�x�,jP����P�����9w�d�tX�ۚ饴0op?#=�m�h�%;��~4�,`s�~"*f��!l��N�Q�Up�~;�7���$ɿa��Y������-��%|�Us�Rc��I�7�Ա��(Ƈ���P�����/p�1/84Y���Q�t�� �g�uF�~h���q ��b'���jdW��Q��t��Y�rQ��z��Hg��f�F�@��s0��h�0G�ڹéV�r�|:)m��.���[\��}�X���C���6��#7A�qZe2���ۨl��g�5��5ߝ�k]J;����� M���Y:fX&~������M�;����Y�c�qۍ��έ�Ϩ�o�G�h���{�����Lv��΀����� n�oS�`A13g����S��Yq��
e(3�ǉ?9�E�Y&���2�n
Q"��p�|�!�7
�N6G��:(���Ͷ�BI� DÅx�� F#�jLa�����L�m�������ɗ>���56��z�m���oc�!�u6n%ǜr�8�?��K7���iA�	e�{��:�b�&�A;C7{�� ��)8'b��S�&i��OM�mKL�S7���t�a�8�מ���9ٝ� �M�ebd�'|��dI��s�@�
ۋ�۬?94�jZlz��� ���qp|ƙ�#1.d����jBY@X��J�Ą7L܁��4��>��Z.
C�?9;��6X���;����!OX����R�W�!\D�c�|i���� 'D�j:w���η��M����M� OO��q����v]��Wn~RȲ_�;�3n��U�wۧ�5���v;M��Ljrb"���J��9���Jj:����b͎'l�+��uP�����y����}����ȑ,y�7��`�v����'�aȐTtf��^ә���`7��w�jq-�	�x�}���S;��b���Y�$�oF�����v��d$����*-�鱸~θ�<��8��H��<����8��4���[�;�Y��pLC�4VY�ڭߦѬFD��sO��6�;gw̑�.LNłs	�X��Ys �1Q�a�т���O����c%�.y0�&�	�� �AC��u> ���(�^Wnth�$�x���SBIU�"�'�sz\V['����ij�9jf6zF�(1iO�z� �	�I�&��!XBf&��/f��IbQ�u��x��M`q]$v'M� Q���r��
�W6u�޵w֔�6���]���A����z�U^� (�3:M�0"o��'m,���3P��hi��\��y�ԙ���q o��o��j2m?���D��~~�t�G^>΄�Lw���Y�VP�5mO�:�s���k=2�Q7��qV��O�8̽+G§����n�{�0�T�-��_��FˤF/�5Y3���g���_���0��%���g@0�K,�g��J/���7t�$ه�5[T��7������d`X��fC��IF��F96�C�  ��49>�Wq�j�i�T|��'��/H����\/\��/����M
(���)��C��a�������\�A9�����bI*61��}���@���a���"'�Q=�N��HB7��Wt���n�MV�X ,4��&cӥ\".���*&��������P�!��h	�"��ԤM�a"{���) Ej��o�:r��
qg��*�%H�@�2Q�e�L��ܵ���Rf!JY���:@#E�Js���+c���X�gP�"H����^�ǅ=#������azm<ޤ2+6�1�����G�)كvkd4x�
���Ĉ�E
�m<�0���J�B�$��g����P��ۛ}u�a,��{{�5*D�3*@�+TB�lJ�=�����H!G�]��������ҌI�C���P@�7sq�;k$�>�s�MȤ�����"	��|�ėG���O�����v:箢+���^� 3��?�:E���y��<OV����1�c�x��Km�q���FQ��qd��8�����a	��N������BCBU3OΖ���+E���� d`�S��'�|k
	���I.m{�CD��1��X!
�.��2�NyA��b%��	!�m�;ڝcV�)��O!���	�6�."�ԉ+Ʒ�2>��*Yf�0��R�-,��EF�&"$ 싑n�px�9)�I�w�yԙhM��2R =�{)�K &�ş{:D'p(w��M#0m40r�����B/$�
&���uD�y�1,�B�N�,�Њá�<"$.���芁V)���u���Y�I�Fa�Τ4��˘k�ʃ}�1�vK�ZE��}�h�
8P��vՓUV�p{�iJ�ϥ�ajv�[�7���u	��\^;��@�(q񿧤�H��垓4��G)� �K�x�����
&�~'�t\�E���P}��Ӊ}�扤$iM���5��:骆��q��U]���I!$���c�b�϶���z����)4��f�Q_iԙ�c����m���z��׶��2&��_��1'( +r�_uyu,D&A$1�S��0A*�N�GC�$���f#P+M�o�J����H��Q��-���F�B{e��H��ěn\YݱԢ!T�Ի�E��4�ɇ .%��耶��d�	k��XY�\B�����	M(s�(;��&l�b��COʙ�$у���l}E�4HVJ��,D5���L�����=4��(rB�3��ax�]�l����	7���}��Ȉn�Lͅ� ñ__ˡ�
��;_wc�4��15��y���$�|t�2���{��]a�e6B� Z8AU�I����賰X�inz��:�V��O��,y��Uu�aQ�$�W���S-����-�s�V0'�.gVu���L�,D9_>�C��n#���-���;�Ue��8XMJ��4� j瘴�#D�`�#s���!\Bi���>� ޢ����N�$N'~��� �k�_��$��//:2O:Os�=߽u>b(;���� ��6J9��ɶ�����K�mI�'�o�$VB�
�!���;�.�Y��2�Daa��N���OQ21����(�@	���������#������4��=@�ۧ���6�������ԁu�z�f��5L�(�mS1�x�@v-]��%ĘRH6��D�<��;�}��@N�>~���s�93Rk���o3���:*�R�& ͱ+q����Ĺk�&53�A�`�������	a�Ƕ�qULM��U��*�;�,n2���KQ�N�lg�� �̳'YË�V�}�����_�Ί��:.>��<H1� ��x�I��T[���=R"s�P�nvޮ/B�L˼��ށ�������D ���j�d�ޱLGq�b�t�d�h�۶2�2h"ZN�7ĵZ���3��my4� $�RY���oF4���,N�Cn�v�؈K�N{�#J�;_�]W����OsK�"$ |g��o]�}���4%L|}�@�u����xo�� �� �\�cC�A��k5:�� ���/^N��B31��0������Զ���t��Tr����j/?z\2���Ӕ� sІ+�"��I�0�Y�}��c@$)�%I��L�&uJ����3��D��&L�G1�[$	g]�/���VO�3�K��u�m��4�L�������$X�8��Veda�yXS��9����uΉ��q�OK��OCs]��nQ�`�f��x'����{���3���$v�xz:@��/y�v��������.f蔽I�t�ɃN��Ǯ��G$ݽ���`LN�K����K������u�b&H����
��9/cl� ��&�� ����ޕ:��o�����AL[�D���tH�,#~*�q�=���T�^}0	ej L��'Z��id�3�U�\�_��j;�(���,��	�ۧ��j^{�=�@@!m�W�]m�	�.k�㶤P��ē�tR��=�/�>��Rrv+����w�}���u[�� ~#�.��zL����gB1Y���i_I�o���"��X;f�mS-�3������1�Oɩ8/\S�Ԧ�O'O�q��tʜ��`����O�ˁė����Vr<��zL�!��D�(��h�o��9���s�j"B��i3�=BUfan�Ckg,��SLH;�mZ�����Մ�-��c���M0��8��_MQTyn<N�L\L��{E̘��ǿ�~ƍ��/N�q��-��H�;׾�6PV@eU��<<�&2�y�S���6��}�t�	��Χ%JLH�����ӂ���7�����PAǟ�+�� $�����zH�+T�o�;����*n�Bح����j��Iy�ڱ� Va�� L��	C�~_ƈ0�q!��o.N�LJ1<'|G&�ht�,�h�Ϳ,�RN[��S@lsGKM�t��lNmRv�e�2[�?�	�L���L1����[��~t�)6�cA0����{���D�2og��a��Lt���i0�D�����oBH�=+�r���d����7��_�}*[��c����H��S����S����>�&��s>1��}ś���ǿ�0�b�Ӏ ��%�����p�� 2��$!9�z��3�x�
�e��V�r`���w�Piy7Б�<�bH����2-��{jz	�\.7��:hQ���M���]�Ƣ�!67�q|j����v����q~�>�gP��;Bq��M�02����$�S�ҘU�N��M�Z�6�2����EL�a#�ѵ�H8����2գ�����E	V)3R�q��3���IeT��Ό�6��������KM(ɑb��9t��a�ͰNf4��u��q�#z�����Q',_�1]w���N���x{JBk3���tG��nX2�n��ϰZK��w._:�KB4�zgЭ ��[E�4�sU�$$u"c�����#�$O��>4�@��s��y � ���o�D��V�L3@8��!דR�#�)"�]�I��G�����6s��A pF�!�3�Aݚp���
 ��0yΞ[�&z��� @�~��}4˕v͝�fu"o�WV~�vl��.����Sd2v5�ǧ}U
�XZ�M���Fɋ� "3[6� ������t�&Ir3���F�����~�f�L�\{5�i���ϑ�D�$�)S�Q7�
E�'�]���"���c�F �T�8�ⴀ�T�P@хl�Τe�˜v���5&��e�����R�u-�,�(UD�t�O�%T �q��1�� Hݙ2�C$� Z���[g��67Љ쓾վ��: uc��j*Ji����^����R%��v�܎�Fjڸ��e�EK	�2�u#��( ��g���$�iD�LS�DJA9����6�����cA���n��_:F%��Q߈��j1e1u�0���Pz(l����&�D��O���@���s�Ƕ�	��\}�G���>��4�%1,T���he��d��gb1�V��2��={^��I�����s+i��fx�� �VX�"Y�N�$ ,b���D�J�m��� ���>#���7}+������S�bf.����J�� �7�>4� �m��� �j3��6v�:�Ξ
F��N�oQv�Fl���D�[�e�g��e�\n�8G��&x
��ϨVF�<$7�\�i�q-#y��CI���z�J f>-�E�G�H�,뽰�z��i"C �<:Z�;�}a1�l��iT���ɗ>f��"D�E�1p�WƦ�w~Y�|u�^�L-��-����4�F��u+:M%��]�4���$3,�4~�A����#��b��a��m�ۈ!D
U���B�@!���̐2g�P#a�g)(�ZD��GG^���.O=�@M� d�4��Ff%3�;��C��F�N/���XĻ"it��U��;89�% �)2,���$���I2&��: Q@��re��{��R�@K$l�4��z�& Yz\��M.����u{�Qow��\[�O�� �f$��M��WI�����N��.ރ�K�#�BK&7�CzcU�D�;~Z�J��fG�k� yCiP��Ɏ��`��V3+Ę�G�Cg(�Eq-�L`AM��W�:x����i&@�%D��{3>5J\�%�m0��%�R��ol�iST��]�y�����y��6':�+`����3�@B�$���ޒ�JU�y&8Ҳ��/�{�-;�&3V��/y'N����3Tv�H�����Ё�+3t��B�52�S��xX	fZ4̩,�n�L�>��Oh�D�L��^�ftI
㬮z�ZP�.Y��}t4������J����r�,����?Ϸ��3�K|h�{F�1'N'ݭ+v����)g57��q�%.�N�A�2+5@���,�⳺i$qC�U�MU]h&��T^}��s� �r�����!����ݘ,���{X�Ǿ���Y�$=O%i�@�5Ԑv{k�d(~5H�Xn#t�4{�!���kҶ��ۿm	� �[��i#)�Q^���2 "�:�x�[�չ��ǟ����"\��|������ ������MD��D�cA@T�ec�I�!��m�]*р�>���˟���5צ��U����p�m�΢�q�ئ8)bH��P!�>cֵfH�8��oK��� �}��o�1��?��� '    !1 AQaq�������� ��  ?�E�/��r��� F�G���~y�+�/�8��d�<��d�L��~{� ���+�~�>��������OK?pN�� �_�ȕ����H���s��|����z���M�6�̰~������n|qV)���O�B?���;�����O��UbXvv���]f��ߕ�p��dྞ����}Y�v���x���E�]�]s�{o��ߞ�}��)�o�ߞz��Y��Pu� ?^O/ԇ� y����b���r���>�꩟��߮R���� \������O��<��_�|��s�>C���k�vx�c���^?'��y���_��;=2���ZC�(�x���� F|pO'�~]�.�x?��c��_��x��T�^��/��9^�����ȶϏ���\���Ǐ��H=��w���[��.�_U��̺��I��<�p�4/�gߕt-�9^����g�+`T3c�'dt�n����/H�H�|�j����Z�f�=�<�>�cO,1�[��j �\�����#b��<��O��&(DwL|r�|�r:)A���@xȇa�'c�x8 Q*[��))�֤q���\k7����{�F�����1@�f,�_\4���B �Eļ:o2DG5�xg��@�����c����OA�o��@��M�oȋ`��!u�L�ƆJf5�*& j+GnW�ڍ����ìe�$C��;Pˤ�Ö�`�.���P��!dT���#5WeU,�7\��U��A2�v�p�㩃#�h�;q��,�2Y4��$E��%�2zf�b!���-\��Lj��HD�	�$����q��n�uo�����7�V]R�� ���"P ���m�.3�f�8��/�9�$UF l3�ϧ h�j�8ҹ�0��
w.���1YUp-f/xp�K��,�2V�߉i�g���@�U�@���0������l��5^�A�0ϓ��0P1|$M�k���H�1�+�x���	L�RL7=~elk���d��5%D`0�>o�g4RO)���3��pL��i:w�ތ`ĩD�=���D �mTE!�p�x�����&7�]�
�- ��W�Fk���n���	���)��Wx><bq�����;8c��D��7���|*��`#��h�D��'"tVӨ"�g�P����d+}��0!Mkِ��KXѢB}�
[@�r�Rl��� �(Jl+��� �c�t\�E�⓹h0I!�eq^#�"��G(��4B@-qJ��F�.#Qy�  ��W T�(C�+���PG4�8J��Ǯp
(v�b�J ,@`Z�Ve��	�ň�D��B$�"5pո`0�`�� ζ���E��fr��[���&Svѫ�`YJ� �͹��Ȉ-��C�%�/�̌DFTn�'E��1�B�r��%����� �r��j�VE��}�n�z]��@s��hPE�|�+���J5Z_�5�9+q;qJ{����qS"�F^O<����ߐ�˩ʅ��n�E�	@x4�[!j�0��������qL)��|l��q!����V�\2�D�-�%6;�N�Ub4P�� �#�fk�KYƬ (�7i\�Ák�v��p-�([�W���z���sƮ4ݷR�*��B�h8 ��%#!�P�i)�������N�.@x�� 9݀h8q0 ��3a�`�M�:&L����L��`�����;h#�ԝ�E��l��VO��6C����׎`ͦ<�_W�1�~[�|���,��i�5��� �_<N� ��<2M&���+���k�F�vx��4|Ђ��Pϊ�\�����TE��8��e�5)�H��D�QG�u��֚�}+��{��Š(Xis}�y�2��)D�����D,��-�q��!D�#���f�J��m��Լ�I���ONB�b�HTY�x��m���(޷&j���d�g#wƔ< }�S���D=��0�0(���!�yB��p_C! c�Rq0���f�:�6�����h4<9Mu�s"�����|^�~�� ����U�HRYT!jf�c� �LeJD�m�q�;2�r�3�3�i"��B��� �E�*aĉ�.7������L�ր��u�uh�E���HӅZ)�؀8���4�"- ��Ȗt̹�p'�ȵ(\D�y&̍�I6����]�t�҅w��x�I	�ޛ���v(V5W!_�8E���Kw��<5��Ϯ���}4S����Q)I�0n���^�80�+�^I ��/῎֔+��p����Q�+���[�0�x	�F�X!_�o*�F�M(�{�����p�HRH�留`+[�\���-���C>N;w��W1	���Eό��7���z˿޵�� I	�J��V��d���Ce�}J-�pJ��A#���I)�����8"S,�L�U��
QK�	P�v�x�D����!xZ�b�*A(��V�$8	O��0�!�0
l'<��!A�rg֞c��ͫ}���塂\5�����5A�g;|��ˡz��|�� �Ĩd7���k��+:L�������g���=y��{�N չ{wN�`$Ojd����N_��Td2��rWu�ѣY�w9�J�M�C��|\���$|RMK SC��N��#C�'� 1��-���h�"Zu���-��g0�P%�	8SP�?t�hR��McI��rU��Z�� 2�TT2�Kښ�K�PQ����/U@�dY��(I0QNl��AK��x���
p�s"����ȳ��L�+�8FW���#Tg
p�be�����+�r6��kfy��$����3̭i�f;{����Uo�u�����vY|����#N�~9��x#��s�a2�~�V�KJ��&���HڷE�LDQ X�-#LrϾ85Q�KѮ$�*P���U`��(�D��>����W#)Ia<�8�2e�QF#J�gz!�8$J�xоH˟��=�̼~O����(Xw={ǮA� �ꥃQ��B��f������".�����<�e]��� |� ��f!����� #�q�g�ࡪ��H�J=R��FTp����䉨��M<gpRJ{[��H;{�<6e3�U�k��<�<'S�����ۋ�:����nn��-%���1��� @69�GƞAm�Q���쾎AFd�b`ޚ0p(
�HS�qw��I�j x�8(9v�D�Y+�]�����U3�s��� ��a��KaLVy�8�Y�(�_8�4zx�OR	�q����e�!���y�W
F��3���d�7��0���`H@Bc@PZ�$������=���Ĳ౐��	��*<Y����0Ai�(��0 0�M�
D��� K�t��`�׎����n�?��E�:�ӟ���Ŭ���x� !��l����n�}'���{Ⲋ�!�kG� 8�*력ߓ���f9�l6f�q9h~�D ߊ�Lg�l��6�Y���*C#++oE
X��I'ּ}u����"ĸ�X���b�����,B����YE��,�R�CTε�����q�5��z՝{�Vʕ!#��Ga��Bˎ�Dآ��.2-�)b4���J#@�I���ʙ���'��>81D�2�˭?�Q|J)�����0F�`-(��S�
7�����p����o��i>��R#���P`�#��C\����}?��Ѷy� ��k<����\��!VG�?N�W�ed�P�B��-s�0����S2�%c|\�b����*�F��ՅŐ�W+�F"�Xx�3�z9�D�K��yhM\�TAq�s���;�Vʑ_���!#e1�H%$��
�(Ȱ�MR��Sf��#*��p@��ki�m"��#�X�/VF8�";�,�V:��tC#���^dG�
�;��`�����{3~ݎ�ďcp%� Tbe�g�K"��` h+}��� V��;���R���n���3��?u�.	8�d��_��&U��f_���_x�>�ʀ��-�"�d�'q
Q���d1�)��l��G���p�jo�5��tW����r]�&f�N���I���
g��a�-�����V#�� �\��$�3{r�]o�4�a���6�_ߓ�U�8��������7�	�`4��M�WQp��/�Lq�+8Y�a�xp+	�g�a#}��E~��� ��������h��"УR�q�+�L�7��ԥ� L�.A��I��z#L�	����_��X�����~� ��+k<�M���$��� �A��}���'���Ϸ�<�vh6���m�#����wŌ+�(�[�Q���խ�T>�X~f?0�/G�Kp�ol\�B�+,�@[�W���@�RS!��[O��@t�s���&��Bj�F� �\�D_)>�JN@�Rp�� ��G=�U��>���}��0B�Z�ȓ\�a`�UCs�e�N$#)��&pa冉��}ȳJ:��\���!�I�7�G�Cex�XFcDS1��ԊܧXx�.>3��#M6G�g���r� _��%VD!}7���{���pS�����*y��������24� o��;yh���0�p�O��C<�g93��1s�N��dϾ�(}��0VhUI \�(U��kj��<��`��G4G;�h�*w��T	�g	�A$��y�]��W�:���
Xj F��y_�@��� �X`���gGc�'x��(����ƚe1�|��D d�Oӗ����0*3k��a*ա�s[1�F��h�� �F؏��n�o�N�I��x��Gw�o��W[��f|?�8���ԝw��;��k�'�C���%�}�ǫ��#�w�?���w_8�yƸ@������x���5�)��u���L2Z��0�/I��+�Yj%�~Itd z����`�Y��2���&�*L,�`�E^A�#A�,�#ae�J����vr�ӓ:a�8J�\�r'6D=�8��Jկ!�j�I aW��"&&�9�,�u�k 2x*6�ܯ��18���'	g\`�E�R�N ��q��D�e9���N�y3TA���E4�!xp�PS G��6�Nq!oo�1��G�0�3���ɱ�O�}x�d����=\m�H�.q��.�.����z��dy)�J���{���C0M|��䘂�A��W��H>�EqJҼ���CZ!&y��D}d���C�C�y�ù�i��;�
��WB����q���`}���'ĵ�pr�  H� ��}�x�0vL�N�z���@@jN��^R��Y�A��n<�c���Q���Y�a.�g1R9v����� ���J ݞ׏�0�j�{�<���'�����L "1�r�����)�2aŗk��o�i&#%}Swf>��nޥ����>���{q���aQ�a6�n����� �um��<-���i��0k&e�b�!����	��~]a��<�H" �Lf�:�9{&>\Cp�Z��T� ��/��
D9[�2�ə���_�s�@�0~��2+*�#ʙf�J��bf��1&�T�E
�-=l��b��5��L*h�xH#�M�5
G�*�$���T !��Rb���� �6�H���xK4{C���*$�cn=��{xEt�-�q�����`���G�.�W��mt;�D�ȟ:�hL+|��rS��
e1���V�
������L���w9�"U���f�̼"S����h`;n�37�ԓ�THV;�7�O\��Ը��ro-"�Y34g��J�\�=�� ���S?(��������H<$��N.�>`X�+&��/��L,��1�sР�oL���C%�����W�����'��<*H/ISP�0�t���`K�9x� @h ��诉_�����ߪ� B�DId����g�IBҧ@T��"��8�=5<G[dH�d�Ù$"v<�j)���
�a�§vK:�ӵ�ģ�^����b�[!���H�<	Q%S B�"z�B--���hJ����qe(\�C[W�r���k)���H�*�JÂZ~���0Ɩ��d��	��5/hsd�.�� 	�M!QE�#Ҧ�@�Z�r� O恜	H��z��MD�e4���M�&H�x�>`_����eb�p��x��D� rQ�1f �<e 8X�{�js~ں��f%��:X��Cef8�Y�ž�LH���W%���*PM"5{7W�-@n�&@���T0\0�M�6�`;w��� +��5��>X3C
����:q3Rm�6����oG3>�%˵&8~��c$YVaN&e$�)�;�)�����w��"$�lc}�=@�FǄ��>9(0ZlU�k��#C��\���8����
1��p��̽E}�H,Ԝِ��a�����#,�%v�W$#_Y��R{�C[��8�������#g�"��eȢ}����� ֵ�0!b,�G���Q�m 3/"wEh�ڕV�FA0��_|T��k���^�^���/��|� ���*��Z����P�ɼf;:�*�Lb��H�Ԡ�H�~S�D�.�C�ۓ�P���o�Љ�T�b9a{%�i��DcL
�b�|�!B��FN�uϧ�*�H�MbM�f�Q�h�Fs4��dQ�:�ߓL�#���Ơ �L� ͇XL�r`�.p�����Xd�J�g�j��M	���\|Y�mb=�����&�2�{���v�HYP����AA�0G�KXx̗���s��1r�!�\��(���J��V(��c`A�go\�es�$!���B�r"�Dþ�>2�X/�2ჿ9���=4'a9�4�x��Zk�+���HC�1 F�9���U2\�ިD�XH�!H�7|�2���z�) I��[N�D�z��r�4tRYn���M�,�2���� ȖY*��X"5�N[J�����!�z�n�rN�8�ǳ���0�+�ǐ�{�ŕX#��Y�Uհ�-i6�=����ٓ����
}��c��H\��{��4hiSX�N����-B�� A00��e���+ D������5Y	����&A�6�S��!��ufϢq�I�.I�cЃƃ@��4
�.�0��pQ����N2
0kD�Pʤ`�X�j!\c�[�_��~��r	Ѐ�0�M=$˹� D���~0Y������m���K�v|<˩$R�����"�qq�kSs⨔)n���~��p�Tzp��Z�E6o�_�7ھ�g����%0��J�'��C+�"�/�\�9K������|~,�As�p2��ο�|qA����ߏ<�x(\}fs;����w���'�\��ϋ.t��n �Qc���u��F8��ߌ>��7A��73�j;ٝ<J 2+������B�U!s�����zC��g�� �~���h�Y_�����໹˿Ǐƈ\S{���� y"��Ǘ?^����"� �ns�H�����q���e�C�ٳGS�¬ݯE�I����G��:>��qa�ߌ�����[�n���y�Ս���^��_����MM�g=���[M���>;�<�q��֩z�ٷ|I��+�}� �x�����4��}� �c���V�z�g�̝W׹��i�Σ��}���g���� N,2�!���޸<ьD��*U���9؛���*�����a���KO��t~�����8XC&�>��qF�m\L��w�(�g"��h{�  �&��^Ǭ�ڿ-�n!��,��x]�r��)�a&xx��Q� ��J�}�[���T��^&��:��g\r\�ܺ�[��uAI����Ӓ;ga<���q;����M���\!�8ξ�@7S�%Vl�����^�Rf��@���NB��n�����K�<Y�N!JYyg��z��'7>Y�?�ԥW��n~���I@lq��ow��Wf��o��O\�6H=�A3��aA3/��ɚ�
�L��g>[덚+�*�TUa��R��폯��Cb_��&��)��Jg~/�́�_���p�+S�񋙎0eps��鯟<N :���ޞH�.[�����P̳"y��n=T�/����8ņ�U�q��0 ��u1��;�������
����C������X:���R�[��療�1���|2���9������s3D������6���c��{�����CL�]M�Uw�� ��t���]z�ʴ�Ҽ�f�Yt��{�RI��0>�ʚ�:.>���^̿>;�O'��S�<��A��N(K�׼���9�[w ��������X���V���S��P�v1Cth�G&v�m[}ߞ	��d��x#B�}��"(�Uu��ƞa�+XPUM�L"���pa!i������HT�9�g�a�����~��$ ��#^�� N�U��V�k�H�>�~�]���zbWM��"��Lj�Ϩ��X�`m�F��:���Ɋ{�:d���q� �JSx߯����B>&j��!���
H�O^��-8�׿�>�!ȟg�o���*I�w���$�Ud.3�7���4�UP�3�� ����fw�?~TJhDc��ݟ�˱y��_�����vs	����3�Z�-��[���w2=h�Gָ���j������E�ޕ=���\\c(.1�q��5c"�߉���yy�"G�U� ��RQ@�/�����O2F><~8TK�u��|CTf�W�ϟ��R,�~>�y�]��^O���
�!��e��.�%�lw�뇈E�B����}���3	�����c������=Nd�Sƻ�<y�x(�1��T,wO���S��M����74�	�_�w�|R�h\�׏����5�S���m6Wn������7�Ưn�6pAPs\�|��s�9Ć�t���hC�A�˿��4����<�����O�� ҟ�7G㿞X�w���p�8�(U���ʕ�fƪ�����U�>_������,�u����@��-�p���L���X&B�ю�2�����8Cm80@��5�TB����<��9�XѠu�5�q��{���殺�c�ן[�N!6ߐ�}k�ĨF�3�n���ƒ5�q� ޸�5<���� P*�5s�M�}�RZF���}w��M.��~��@�g�� ���y��aY`������˧Sپ{ͨ�}z��ï�2z��,�޷����Jpm7h����(8o_׉�d�=�����yD�I���\�Bgӂ=y��9$T.N�,+��$y���u� �
�=ya�Oƹ�Ŏ�Xq��8a-	�A��k��CZ��X�
�~�����s�~=�_1Z���>����@��w��<|r�K.uO���)B����P@3��hȸ��: ���^��� a������Ϋ��SD�X�!����n��?E:�|I<�Q�L�8����2��߬�?:d�=�����G����@^d�~�M~���@_���L��@B�ƭ�՞9H%+c�3��x��P�?�q�*etۗ� �A��ž_�� 2}q� vp�R���f�bq���0�c�g��&+ӝ�����"������1r�����	REi�J�y���X�@u�,	 #PU�?�`-QP��W4'.�����|rD��h8����3�U�ku�美A�PP� /�\1bc��eQ���r2X������Փ"-bB�i��BAD�%у�x^`D��wۋ��dLgO�W9��Zc�:�:��ښ2��a?���c�j�`nD ���-��Љ �4d�^4[�}-8@� 3��yш}x��D��)��=��#���X�Y>�^6|���0�y�/������)׋�J	*�QW���<�0����� >�hJ��F��xU �5������3qY��>Ϡ�1CQ\��G��*ͧ�����5>j���<��=μ:�ϑG5��94?��uF�
v��_;���J�pw��⥕��u�~y�L��t�7��]� ��.Q�r��D] -k!*�l]w�����[�2(CY(�J��Dq
X2�2�W~��P�:�a2(� (r��d3�GH ��B�� ����9~�ڈј�!�-��4�l���Er�w��i�"���2�z�듯s���LF\���b0O���|9�a�?�?�Ę�2f|}�tռf�P�N�R=1����R�"#Zc��3L�E��r�o����mu[�u�5���a�����z#��H0wk3x���]܌�^,�r	a3�(qH�0�ש�!�Ms��u�<]�&����3�cDt7o�wI��LQ�湳_�xT��<�)�;�mrr��m0de��n�{܋ycͨ��`cb�ŗD�iD�N`OJSZ�@�q8,i���/���;3�!������%�ZA�xФ��X�	���CP�[�{�ĺ�0��;�~u�a�U�s�噁��L�_�'�lB�N{�}Py:[K]{�2�mn�޶���1�1ß���"��Eߎ?�+�珚����~�lK߳_�`������Ǣ�2���_���V�ǩ�ׯ<�FN��g��x�KW��V��_�\m����<r�W̾�y�k�Is�j&F��'�!'m2Q�>=�D	P ��<����n~B�,DH�0[�[���u�g�N��R�!�
�9���x��1���#:k�Je D $k�K��}�Ppeц![�
l^ˊ�1�L��d5�n���&�������&3Ҩ���B��1��:����=q����O�9P��a��L{�F`��A\�<#�F"Fr ��kO|��C��DL��O>��"1qXDq;�8eL*�dC��q����_�I�"I	%`�fz�;�ݶ�_n�`���e��Az��3������Ӭ�e՜�L�����ϗ�lPL�BBhb��1�D��\G<�N2҃ɓ���k�_�YM|�H1�y� B����5��� ��7Iѹ����FaQ%�/i���)�4����4�)u�\xs�Rdz�� 2�d�"��V��ߘE۔'M}��$�O�T`J�hf��������n[a���!�s���略�G=�n[�|X-��\x��\ߪ�;��#|�\zÎ&gt�Ç{O�qQbuI��yFd�x�->���	������S4�6�^={�1X3�|}!��c:����p`�piA2GZc%��׃� c,8B���B�3�P�UU�)�_A��j\^��  *$�5��z�(�d�pϰNLP*MH_�ěՎQ6��;�%���U� k	^�im|~8.���\ �8���D`𱳗�f�����F#Sd��V��V�0��<D�!�A�_��9
��ﯮxJe|
�t�j�8�� ������$��8-mb�>��?�� 9J��s|g�^P�iX@з8p�,V�#bnk�{r�X��<}�f�x>0��=����@��T�w_����?�v�||m�����Ə��˫��:�� �YcD(�p7NkC�4�jMA�~�ؠ@Ʒ���d0Nc�k��"����/v����{|�D��aS�����.�#!	Z�^]~� n�<�B�e���ŀS,FUǩoz�Y[�����Y�I��p�C�^cK���?���C�|��w�>�~>��4O�=�l���8r��w��� ��>_���u�"Ի身q����{��᠄7��}/[�� @��>�^(͆�|��9d�����䡸[I��|u8�+�U;� �� N������p�U�7wY��Q֖�}fX���G�gɡ	�@�e��F�Vc��Zaq����jd �Lj-�¹~�A`u�5����r9������Mb�*�I�%�n���.y��%9��m|�A)���A2���8�˹�	R��ead��M�E�p��0ԝ�a�٢kI�.[��|,(a�� _|qUBV� �و�y@3XQ��^��"h�x�
��#�3%�T�������������E�q�zz��(s���I��B�1��D`�L��
�p�Fc����!����w̪ ����<E(�3��~|q�0�n�+w�_OvcJ�����0[1RЇ!���I�8E0V-�:&7�Q�iڕ�3BWN]��rj��gh ��o��(�SƼ�BO#�v�.f�ɛ�~��0���ՊuH���R�3�jM�2�;���18Q[d[���E8l�P�G偓}h�B0�	��o�+\i���N�� 9d�6I�-R��*��]v�qT��f_o������|.\��Ipb�[)����m���:�ќ��ߏ�Z ��;���/"c��:\��/(�a`޽`����펻�?~Ggo�q��dt[�L�Æ�B
&�;���1Cý�ޱ�|[�H�De煃��d>��#�4(!t��Ŀ;��!�P����CWEEV#�R�â���� �d��i�B�;�%�@�4�Š��S!���Yb�֊BH4C1����f���x˭�qZ*3)�l^YO(*�gq�!���<���ן��bj�{��7�_���),�2�� ���"�Q����Ɉ�N��ӕ@C#S���s������A����г8,�� \J������w��R��LR3|���bw	� i�)j(�I�E�7��=gf�w~��ù敽~�7�ٝo��ⶋ�>]>�n^�&�9S���P��e� lP���'|��D�6�}c�xJ�@���e��k��A���ξ)0v�f�i� �W�N��^���_ �z�w��}���Âh3&q��
�e�����"�
�� �y��1��%�{�c�SG�SKr�Pڛ{�pR k��Kc4o��mΫ��?� F�חx��p�W����3�u�p9����q�8�7W����9Ըq��y,�D�������]���3�٘{=��e�F�zs7���JZ��S~�*@M?��h�����_��e۟��Q;~��z�plǽe=}��	h2ri;���.�Ǚ�k�}qA!X`)Z
��=yD�D���׮EHdX���O1�":�I�����p�F�n�7�k��l^V0�ɣ�����r��?^�bV��}�q��I�7�`~7�B ����iz�!�A�g����@Dӏ?�@��OWo׮1$� ��ht8��Y����>��Y\U��� /�"�W	�� \�0��<-1���N黑� ��&��XZO~O��z���U�|�MUl@��p�x��=�(�$ʊ��/M ��0��=���gհ)���	Vk�u��	f���Y���d ;�VX�ǎF"�xI��]������x��Ʈ_��pgo� 8V�j)�C�}�� Ѵ*��'F�AƖZ���?�@��$&�f��r�I��=\n'P V�a���J��"
"�P�w�M¦꼏D�m��h��g��	Q�n��__�+;
mX�a�=�{��e���>�yt���������p�V��:��
�L�S��<w��0�����x�ȟW�w����")����ƍw�x�,�<C~��qD�Aq�o�_�Kr�����j	;k�/�(]����Y�#�A��q����||kX<w��I�I���g^8��R��o��)t�>	���|�\[����p����L�z�Q	������ <L$�����ASX\qRE���H@g]��ʓ��tw3ªCԯ�� ?���Gb�.u��e�3���� |rd����3+�x6W��1j	���2����� i�T�	Ly��h��� a�~v�O�"0�߉��n���7������*5#߀㌒�H��'	��È�T�1��X.r-l�~�N/+Ȫ�1'h�/	�S*�:�
����.-|��4#�����] �� 2����I2V�����������ịV������Q�y7.&�/��f����X�b�򓹎`2z;�v��.jCH�w'%�*P"���Ļ�[z�>�;G'�"�
�*A�Cu��BC���t,U��|Dl�q�"�'������IW���iAf��iw�L� Z��������eV-�fK�:��5s$�,�[a��)�w� 9�&pm������o?�:��P����s���0�I���*�<��_��ɢӌb~�E\���?q�Pٯe��n�,�<�:�sg��9ˮ,Y0�a�ǃƸ�z�~=���g~���Y��_>�C������ �0�$���҃� _���� k�� �sA������B��1�nq�q(�N0�a�c����ܕ�7��ӄ��y0
x/��WTݖ�)�s��dL;����:/����}�9hL����X���J�-R��%U��m�g\p8����c�|^V哸?�Ɠ�[����1Յ2K�gz?>8���}����)��H9ApBϯsQ�!�QFEɛ�j}D蹏�ߪ��dXO;��d!\���>��ɹ�CJ�./�� 0�ԕG}rB%5�db�����=�&U�x��b��Q 	�8 bpYtE��֋�v�"hk�"�鹿�:�b�`�@��Ʈ;��� {q<B��(�u��� �:��Pq��]`��{u��?�.6���v���5ju�?f8q:��c����>|g�
�Z�k�?^S.}P9ű��T�+��� .d����ɾ \9A�?<bF�\4��'��VP��� i:����g\^�t=~�_�fl� ܘ�u� þ�\E��>7� 9�3�������xi��l������'�Pam�D��2�w�V{�� �Q�3����t�%1�.�ߟ�W ��v��|4��4.�0
�i��~>6r���w��Sp˦g�<P�
Y�t����d1
u�B�����`�G9:�A���K�8f>x�c6k�z��&(����{�-o�e�����>�i�;��AL>Y�d���+�Z�� `��!,�:Ͼ.)܇~���0`�Ȁ�p1�e�(�ޥuH b�,m^kN�N��a,
�c�_�ya�dF�i	��\�_��֕Ԩu�Ov�P��Z�k��df�� ���� �ۮP
m|�7�^�y%���޳8���K��� �\�G\T{ߍw�k����ߋ�|�NŲ�}y�%�D��I�(������ 
��>��8-Xu�����qG�~w�������c�x���/��������^e\����)g��0����!�w2�c?���??����d����c��mP��֟�(������}q�c$���j'W��� �����G߅��\�,<ɷ�^ oD`�f1���U@��!rN2˰5�s̻?'��ۙ)\��&���BEq�$�pv��e�	zR��yᰬ;�����H)Y߭���/�ˬã:}p�n\zͿ�y(L������(���k�y:f� ��z�ĢG�5�'ӎ(�a�s����o�!H���'�C�O;��I{��UA�0�a�.��	�p�X�4;=]�j� ^@��! �886rCjRM7�q�*LN�vA��|���Me�QRHD@�|e��7�[��l�)Sj�ي"� L1�Q_搐�Fh�@�����B�Ԝ�}ٖ��Μ'|^P��Iӝ��r⩠�oD6���kʝ�^n��U͸��x�C�S�����1M���B�cߛ����\~f/����g��}z��E����~?O�"�d�\w� �1߃����Zq�� �MS�\ ��?�댌b'�Y�� �"�8��W�}s& ?_�?kF\}�_5����<�1�k4�5��?�|eZ%�D3<��$�� ���qf�f��#N� �z�S��;%��?o$������q��6�*����Xv����<M,�|�AP Va�;SH�z�ߛy-f�fg�?�9�$��ߟ�&�wݽ�~2k�MW;�~���4]���R�� ϊc�>�.��v�-F� YNP&��A) #�d�0@Oj�Z!h�����`�C����P�(�Ӏ1�`�"�l�̅@%-��,g����9�ҹy$�
��U�Vr}5!:A,��zP̽|�p��OfCi�*�`em����M�Eg�Y4)2���e�@V+�|�XJQhͅa^K��m�iq�P=�L�f6���V3��E��]���\�=��dZ3�e�Rt�Z�TA̯QD�>�8�C���y
��	BL�b�E�M��a�>��1��W�x��sf,��c��9R�ߺ�Y��\Y���qT�Q+>����@����|p���N�C"� ��`+Y�m�5��� �|{��� ���@�]:�����Ϝ�#�z�����
���z�@���a�����``�c�� �*�����J���7�rq"��o�q�H!у��� �x!�����110d�^	��!��Q��}]q(��4���P��4Y��5��R���X��ι0�{a0��� ��`��[�+����63��h�s9,Y#��}�u�t�y��ɨޗ�}|~�")��n'�ǜ�DÁ��b����7e,ku�_���i�@���A�Ky~y�6�fG�Nj6J�Xy��{��XBA��7 �,P�2z��	���S��uuH4��}�ڭ����;*�$rƃTb��L�6�M<�G[IIZ9R���ST����+�\�;Q�����t!�7�Z}��KL hs��j�p�#�'
��E��1������+Zڊ\X�׭N1楲-�3D	���.C���Q���f��C�ND.x�h,N��8��ؚr�'Z��-����V;�
8��N�
'�\S�(Z!@1rDM��ȌV��B��w���p̪�xB�Ƿ��x�o�)U�E����w�s#��2e�vr�f�����LG�����6&�M�pEBV������ׄԨ� l�zwő��!��J�,pJ��2��wƄB4������
�� ������s�1����1�	������;��N�z�˼A&
m��4~x�-n��w�C�@~��r��� �Ĭ���+
��|��f"�iL���2A&�LCG��`B��UK��j�65mV���?�W$�5����G0���\u�	F������h�s]>/fx���O�y?^Lec��yː�6����ł���nr�˨X
q7��bc�F�q�{Ã�B����
�����:~�ۋ�O�P�4n�+Ʋp�k�nd
ߍ�Q�fp#]�C�1�(������1����jT(���ʈ���ڥev�
���I�	�V�
���� ���h�"`l<W ����`cy��H D�b<��H	�p�����H�e}���(%0�6��X<N�R�$� �e���0pT�(^�_b�l�*#\M�"~�����P25�Ԫ�jW<���>� ��0Rq����im���bP��+u������k8P2�ًrx+K|���PZ�����P��x�Jqzdp&^a��$�C�����:E��GsXҕt}�!r����֮'�X�����L���b$n������"����Z����ޱ��~9�4�zO����+XcYo�9��5�a��Φ]� | �"�ł��{�|�t��l
,�b��ak��r K�O/�@�{��??��r!T�%�S-2�J�X)�fXV�q elC�f!���dD��h�Y�H�1�/_|��twxө�� �\ۄ�v`U���
�����r��5G�B2��g�;�N)�\�&7�����R}��;���GRb�@����0	� T ��Q�f�Ǒǿ��)��X�8�� �T,C�6M�x?{[x��#�M�(�Q7 �G�Ӓ�1�~`柄�@$��{{��D+�`j�'؈6�4�8� h�2�2�@���鬅)�^6�9$�N��}���YXTV�pF�N@��N�1	xђ�-�Pқ�k��%�抬m	H"Y�XU���k���,�.1J/�'na����#��h�
�l��4�1.*���p�#J%g�8F��
��Ӭ��Ȼ�DdⰦ�j��,JqYy
�VBG��"�A�1e��+ �P�QJ1|��.� "b�,:� �0C���4�
Pm����獦��+���4���r��$ � >p�
	ȭc(� @�{�;0���@�b�-<?�G2��ۏ��� sd:u��R� #-|c&��� �	�8�z���E ��	���XȊ�u �y�2� +�1�x�1�~�� \����)P��th�����}C@QHv�یrD�TT�=3:@jڬIU�S�w9Pڤ���'�9!EAq�o� 3��;"�:���&�� H���㊕���%.:=�9��ł��ӈ�"�I�u��Uw���e��\��/�3"���I����3i���Ƀ�oY��9�*��w_�e�X�-��S���/e%���u/~���Zt�~<��s0\(e��|q�X3�,��9;�.x-����S�]p�L�p`o5@�y>bŁ�5`�aEd��)�I�#�$0�
Q|J�l"���nr�8ԦF��=�ᑃo�)^���O\��,ҠY�q_(Z]�d:�/�Y���tB��}rT���D��І�9�DLH /��V	��$/GLS�j ?0�X&5�f�JTP�Z�� h�r�7?W�43�o���@���o�j�x~L��P�L��>8�¡$s���o#Ƥpl<����u/Ǟ���c���q9���>����l/��5�+�8��� �9P\-���0��P�� �����k����� �����$�~N:���"}���6�Ah$h�.O<L}�������x*"Q\I���C?��*8y��À DC���dp�B'Q֔F9s8!�l��Q����D�]>\}�����1���|r} �1O��4cw&_���E#�>?�̄q�C�x����]��.&O�����]�u�p)-�;��W���]xv�o�iJ����V^JR�3u���]�''c�8�iη�b���_�^�?Y����Q�	���rH� �W�}�sǳ�Ș"C2S�.�D�m��r��� wAn����Nd�D8�\f�
ˆFsʧM�$��|�� �AE<��(M`xh@�M�`&{HѶ�o
b+�&��T��r-��G�=p͢�/=��j��ֈ�3��+���v��A!G
��'��uQ8"D�"=Y�"x���T�6����D�+Q�<�'�?7�� �=7�@!���(L4�9?����=���,�� :��������6����C�&����[HN���}� �p
��ǿ��tS����ݯ���A2�49��O��$V�%SBt=NE�|��<)dn(A�����!@ :T�IR�ʚ�P�K^���||�y��!�2�z���xu�X)�_=f�>lW����.=�De��m>�'�@����d���� rd�� �o���4h]g6e��<��3��4�9DI�k��~g1ś���.���(DM!��^��0T�4s���[s����^�a������p�jk���3΋������-f�y�5E
2S�O%�$�ѣ"h�3�1��4b�ɲ)cd���g�ɶĮ/Mc��q%.�ԨelZ` �pK�皞-�F�0"��Z��q��̤ ��O�P�f`�p3��`�x������e�~��B��W!(������jpj~FHØ8��њ�xQ3��| `xW�  Pb� <���t��
Fʿ_G���������'-xw�o�$��ɢ�f=�&�0ZY���5���Ve�Õ"ɘ����%.s8	����߆��%�����B�ɱ=H�䒣]�de�G�|e�@��(��d���v�H��T�*zQ�������e
3-�. �!�3�q�A2�cZ��x������1ê��_� �2�h:�&�I�����˨���>�Zx�'h��+M����t�ν�Ւ�	�����S����x�D5_�����'��?�|���
�0��>9��~q�_�1B�S��"���Y�� _9�+�R����
�]�|>@�"�il� y���(4��Ǜ��(���	��{/3H S�r�D�b��!^vciؔ�N5<�G=�#��o�`6�9��dE	�865�V�e5QH�K�,����u��7����g�J�#�)A�)��ܔ�,!H�OI/L9p�*���`� %y�"��&);��4p�,!��*R�
�R�.� �۞%[\|� _��E( �����Y���Du��� >��tvj_������
�<w�G,Du�I-E��?��BSV|����H� Ҟ�+�<2B4�4�Z"x#���A/I.��d������u�����X]�bq��Ÿ0Xf;0U-AU�!���)�'YUk�W?�%��<�����I>|�rg��t�k��Y�-�-�~|���MCx�g��� 2n-ǯ^?0|}S�ǮEV��>��U �ߙ� 1�XL��>[�p�ML�ы)������ߊBN��=���*�;��=�d���ݓW��ޓ��w?�r����=q��#1�1�>��W���ɟ�.��#��>x;B����W��u�1Y����*���}I�3Ȝ�)4��p(M�S������?�*$/Y�=���� �/�L�q�Ʉ�2+�V��9}Vb�S����x��̬S1�M�� x������Q �.b�ޒ�q�hG�������M��Y�B&0�e� ���"
)�~s=N�@�����_���J6|�/���
�������~I�8�x��w�� �� 44�Ps����z�}\�Q;�j���5�1?D>Ɵ}}�@B_~�>z� ,vFy糙2Pk��g� ).B?��ߏ�DIQ������z(a*�XrugQu�z`g�T4M>	�{��t9}<!�(b�B���58w�)L����a ����T�e3�}>�M��X�9f	&q�{'���N����r|~>�0M*#'bm֜~堍��u{�� �Ǔ�:��_�T�~�O��F�p:i�U��8�԰�D���!LQ �Z]���l�,r�"�L� �q�����=�P< ��ٴ}�<`�,Wl������w�����Y:�����*�#�~��?�b�h�qYMc�:>��8�P��6��k[����\4C>���gÁ��e��k�qP=h�U�m/!��67J$B��iA��)+��77��J��D�V	Z��&Ÿ���{�=�u�"/�=μp�8Q�X����	@�����L�Uj�o.?���m�w���AZ[-��?�z:�,�A����������L�t�"sgׂf �B�^5������P/(>�f�cp�p�<��S��pB���!�&�+�@pm��g����,C�xu8�O\��0��Vk�PژN���r�0�!�T�{`a.���&�1�^� ���)uO\��o������@
��� s�0
@b��3� �X7N�rV���}��pz����`�G���ёq8�a��E.�Tx��ᯅ�M��xA�&�9:~�e�sB8ќ�ׅ��g.?�����E���Y�z��F�E��{ �p�� ~�|�Hr���.��x�L��f^(V�"ْ�؅�y t�� 䇹�#�*��4"J L
���w�H5��8Z7J⢛�J�^��I����O���{� �� Po�A�� �K�23:��}e����;ܾ���s\���r8�o����rs�8�©���j�DR�`!2�]�86�ZB. ��1S)n/�b�a��.<g��d;MU��\�6xN���� �E����2c��$?��������"G�<Y>A�{�2�� ��q�~q������O%UI��3G��J�A�X#��_?� j��XP	��T�;5>@�rK��`6a9@	�'�6�r�D8VZa�� {��@�f��%�U@L -Ǧ0L|�$&s�|� =��{}���Ӭ��?'�afT7�G��B�y�-�%Σ����2�@�����?7��}���K@IIC03>���o�Vyse���k�E����B�䣓��;����n?�ӱ�u�1� �8&��._S�{�xû[�����9z.J� ��?y6C,+��~���*�V( ���V�YUGD �0��TH ��b��P-���G\�<�����-\��$<e "-	�!��jpEG[� �t�?<��?�\_W�@������`��1\?� +�k���)�߯��e�c�T��|B��xo*F��T2  Y��(,'Br�Z6R&A\���'�b�4��Q�o�� g�o!\�����{� �� )Q��Uj���#�)4L�W��r�Z�$����vj��$�P�8T�������u[�0�[bIx/�*
���@P�h�i�M�"ł���^ I�{�R�'i�hsPr*;�p�����z�LZ��	k������ xF���.��N(��+Ooxx���!��υ�8����>ЀЩ�x��̮߷��r���w�V2;1@�o������P�!�r:2�#��֞"�3ϧ����*ׅ��[����?���X�g/���q��B��}���n�M�9�ߎ*�"Y�y�c|#b��
PA2�YmT�%B��,���� 
P�.:5`Zdk\�T�R�}nK��y�/PЅJ�Ez c���&+.��g�ZǓC�� �E��ر���熲�ȕs�� ��������5�\�16�� �@b�l>oߎ*k731�X�W�x��b1��<*�1�L
G$Ǥ�~� ��p(,��b%��;�Ry8��~u�'��Uk� �ˮ��?;�� �L����}?�k�1`����!�t@XA���`��A*I��3�J�.��vXTm���M:vR�D]��Ԟ��e��rr���ldL��YI��/�ᑬjQ�g�Z\�@ 4P.M �=w,-�z;��pb>�[�x3���,H�}��:��ſAp1���Z��h�4i�rW���;�1����$�nC�p�OW3�e�� ʊ�T�8�����X�xɟ}�菪�r�5�(P�ط;�r�w�|�q(�9�Y�վ��B�U�����0��a���cλ�W��=o��ƑDW'pk�s����jʸ�OB�,A�W;c %4Q	Xkg��
�T�0��w�D��/�v��nCh0���~8�����~����>�� ��*� �����=s����ξ�?� `K�q��rTDq?~�'��Ҙ�l����$43g�q��"Ү Hq�fE(b$!�ǠsC xb'���N
�3�|�r�dǯ?]��?��)PT�~�%��6� W��� �-�W� 62��� }pڊ�C��N��� I�Hv圭V{��wn�4�;�b�������-#�*n ��0 �/ ���w�p.�c���.+&�J��#F+��' ��g��s��L�u����E�n
g7��º �#߷��C4NIF\�o���(7L!/��k����vK���@`�섣b`�� ��D�^[eLk�aφd�tU�p���l�Lu�r��T��3+�� 7�񾸨���S���� k�	���w�"|a�4�o׍�X��>\�/�����X�0x��������z��f��)LK:ǖߛ�d����_��*D4�b����^D����ǯ� C�/�﫠�)U�K-֩���ǿ��ND�S:?�'��K���>�� ;gv_�*���,=� �pA��^,��{@����=���s��ۿ�0D\��,a�
C���u��[��_(/�����,��s޹�".q��c��<-R㫽/� x����ғ��&���{���YC���W������x<�a���������>:�{�Ğ�}��6��/��r�J����v��������A���~���������ƛ!��Az����+5D��3=���1�}S�,�6	ӳ{�� s� NeU�n��׮P����qU����?�J�kK�g��p�+y�Q������*���z���x�Q*aK&q�!������� V�g7����/	
��Z�\d��P�\��e\��|^��9Gd�c����q�@�����gņ>��UVTR����4��刧*C@D+�..b���ɗ&��5Âq����u��(�6��������{Pi��q���x5�̝�@�ׂ{�=g�Ȥ��*���VW�&��x,F�t�Χ  "ƣ��8&���9g�"���G� ���ҳ�� ~� ��寬'���)H�o���K1s֟>w| �*�qOϧ���"�o���LWG�m����L��Vx�K�4�u�f�l�� oS�ߛ���+hӻ�C��� nj�/�^�|�@q.��L?�W��͜��!N��v��	c��{�u�߿m�U��ᛛ�p��ǽx4��2����lüm��d��2x����$�`�O}��"홾~�SYT��e���qpm��/~5D׊ߜ���[��=x�fT�����!P�w���<8 �/���Ƃ��e�;��s�Z�ɕ��G�Y���@2|��� ��'
d�i~el�Ә�3��&3����2ۅ��|q�i����
���_��z,���ZD�g� 8x/�_W_~�%L�H�l\Xm���₾G.��D<�A�}Wc����|�� �2�g/��x�P���U�2i珑��M��b�9w1Cf�\�1�l7:v�s��Pt00����\}� }`kR�|�9]����s��8��WF8A	K�k���N�+��W����n~1��I�x2c����9���� 3�z�3�E=� ׎
e�E����A�|~�(c�� s���'�=<�[�� 8)d
�u�Q�8#D��L���� ģ'��:�
b�>��~8�֋�����L'�~� |�8r ��*n����g7���7�/�3��L=ۯ��8��G#��%�~z׍��<�3q���٫�z�. [�G�.�����p��� \�#�N���pa8i;���� �����:��'���J..O�r�f����'ZW.[����ķ%^�x���8GK��m�K��?}pD����_8 �c�.{��qB)�������	�r�R��7�����J�z�~�������re|�����
!������\�d��w��`9�J��-S�y�(��sMaRvh��Y���� �� ��J�I������znɪ.�����e�2g�J�
\�)tyK�ʅ�"Ua|Պ��mҍ�Q
3���qIPЩ�8t�Y6fG}Hz�A!m�f��o�����h�� ��&|�8�̰��s�՜�����*�w��G\'#cG{	�,�$����1@���NR�~�-"�7�
ܛ��(@���]�8�i*�Cx��I��y5�g��ۡJ��9��A�)��)d�s��gQ��#@��w��+8cY�V8��x�@��o�����i� �����?S����6 y���mr,=V��x;��ξ6}Vp��Jj� ��i���KX\}���U��|J9��0"���g�O��='�������ZTδ�$��pҪտ�_n����A���wp/!l�;��|q!02��iY�<lZ�=m��|���pũ���P���1����1��?n U�:n]~������ ��AH���\p�*0���Y��&|r� ƂZ,wϧ���Q_EsF��я���C����㒨`.�|�oϸMc���6�>9G�Y��Ez����-��_0+4��^�N�3mU~� �¿����}����WT�1�Yi�9�������F,�$�S��"�;��J�5�B���CD=(�}g���`8�w/-����BQ��uN$QJ�w��+���9mڹ�O(�)8B��bE�gY!1�\,a`�C2�q�E�I.Hf2g�Rhd VM�	�����
b�q��0��.V�x�e�R	�tϿxN1*bL`w8�bY�"b��e�x� @ ��!N<�fB�rj�� 
��(��	���5�Dj�p(B�%(�(�	����Xe9�z�]�9T�W�w�)b�Y%]pR�J3;1m	�3���8�T��)�K�������J�o�
��rs�U�A�kN�0/b��N�O"�����WW�	�U�m}�!�f564&�����JX@#1%K� P`�	H�W9���K#3,f�@�A�K2�	N���X&PM��� bL���_#�`:
"jY���&,ݒZ�q4�(�H�>E�y�X�W5�r���,8�f�N?M��t�:NUDme��g�����&�Ăl{�#N���?r$�M���-���	d�N�|*��s��
��W�D����.���0��a��l�>�b��j��D ܜm_f|������/,�FׂA%�F�'��nRЇK9�賫g��z�ˉ��xHLP0L=��Mp��P#r�bfk�W��`_�r�4R��E:�qp`sg[bJ)�\ZF����~�����Ӄj�����p��@ǰN�x/�N�Y�a	/[$��J�\r���ATm(N g*�� >�`F�,�k2�/�C�,i'���P�)3t�i�� �!ˆ�
�A�Is:�NbEaUF �JP[�8�@�^3}�5���1�y|NAT��L� �Q��\Â��S���"Vi��Q��$�
��@�x֙x '*�z�$6��WC���U�1�<54��)si%��Lb��E�;�8��U�c ���ݤ"��L8����,�sm�����D�ࠅ�Q��,�ޙ!�����s`DQ���%�=��s n�r��b1cʎr�I �>̫s#�D&`[�w��`q-h�8�q�FS" .���c�FYi4������{�=�6̼1	"D\��i��s��C�j�8^�*��c�%�Z��9�\^� /T��K=u��҄Օ�T%2�Fw�h�B�/��dKL�N���&40��|i��\�)�z^��B��T$*+:�e�V�)�*{�hQ���5�c5@�Jh����P��Gf���y��i~��X���]J��]���Q�"�r-��[���Jx.h�Dl8���
��g��Z7&���/!��N�P�c<��g{�������-���� �w���b�Y�׀��xc@4i�\z�*yC��^xL�^'G�񇂸��|Z�pG�,`0�c�o��$�A�<���i���#��*�U����4.2?��c�<x��u��YHҍ�\tָF�Fɋ}��G�X1��=�ώ����y���!ÌuDB�Xy���J�'���,�/m��{y���t�iW�ٜ�6�a1��k����F`�{']�Q�G/f��l/r�r0d���`]��(��x)2d�&C8��p"�yɘ7ܐ��� �(2hP�w�"(C���pf�,*rB�|o�{R���WZ&@�Ţ�X]ه*��V�e��ă�rk�v� ����,
2�!sfx"E�aF�ߏ�	Rv��-�������d��c�q]L�̆n�>8������;48~uKCL�����	��6�1�5�|y}mRA���[[�PH{X8�F��|�>#L ���s�rJ�4�׻���"P>5��&����/�
�d���G�)��u��Z�J�2-�t��|��']r�a�0rp�rc��6>����
��/�8�T�rT҂�9� ��3�7�r{�4.3:1��'�Dsm��0�c�� 1���}g<��7W�O��|)3l��]<��;D �3�
T�hz�:���ʬC�Rc$�#�������ܼl��|�z� I#3���h�%�P�Ŵ�4���š/!�y߿�ڬl,�����%	pp�g�g	3ϴi�	��3&��Ҫ=4x���]�H�3�� ���w?ҁ.T�#>Q���q�b���}c����'$����I2n+��	�߯�5;��Vy�؍��+����5$i���� �-hf_Q?m 4�e�<w�rU.he��7��'G����im���A4%���A���5x�1�9�=��0�w={ケ�����cQ�2�P�����k0�ؤ�����g�a)^��N T��GQ���:�QH���I���"d䞃�19�:��Ծf�U��0�~�����"S(��9ok#���M�$����>�8��]���ϯ��/��׉,� x�ann��|�d�F�.BR��b@��L�vp�����<��>��'�61�*�\v-iV��@JΨ0��u� ���L�7�xJqA�tzz��lXrvudo�N+����_}wǁ���lu�MJk��\�� ٮ �ls��瀄�,�+_Fqb ���}���#����A!�J 7����$Wf��H�db	�����N�Ql�C�|��#]����\�T��'��|s��Sws�
D�����NdU�T�������9��0_p*@V�;�����+3��<��\Ld�t�
��ժ��D�߄S��i`L�[�5�2P4O��Wy�GT�is�4jQr�_��EA1
&*�C�η!OD�A�r�q��l��&n8�R�
ђh��] ��p�z��L�a9�ӯz�H��D
�e�|k�Kr�qM�����!��:�����'�rI�hQ�Zf:㣱3�q._fC�J�O�8�2���}��"e$�b;~� �`�A�(5#��8u�#YF�=5�d̹��:���t���7����6�QL���(�?� `C9��z ]^�� 2��z���|{;�=z����e�??u8\�B�6A��5��+%�^ ��陞��\s=�8Q87�	p�߸�-�P��I9n����9��/A��:+�^'��A���C��F�54��(�>�GlΠ��l	����i#��.'!\?�~�}���0&�~��HCȶV��+k�,P�a�n�"7�@�ȝ�����qXQDTW0��`�Yz���X��0Xkkxt���2o��TZ�ͷ֣����0��=�u���S	�g���t@�S;�˭|r`�&=���ct�&F�.���<I4�Sa^A��s#�% .����.�b��*�� mAJ�+.>3������ӊ�p8)6r$Q�n�������AꇾP�GJ����O�9`H�/f��� ��*����Iz�������r�1	�/�~<�)L���9�e���o��㍚J�ҽ�߽�V��$��^�;��0�R�F���V�/y���B���*�=���4�H¿l��_G��pه�x(��/��㈘�y�� ����?Q���8�+��P��{�?��t��hꝣFrC E`,iwM�ȁ��Ɍ�o���>�;��|��\
2����n]��c���o���0�Yt�_��*��AuQ��I�AU�X�A�i`N�����w��~����E\�ь�%��u�j#P��B "�Y�1A�)���S>�g�vѤD��LsfE�^'2x5x!����ޯ(-��8Tuc`���Ɵ��I��[E�|� x9�&�m\i�1�ʤ ��P�e��90�Q�����D�Y��v�Y��1�V�Մ���6g֫<K�*%���u����񮋂d�f:�3��X'Yv��s$��ڊ���_熓Ze����u17�^�$��y�`�t������j�:OL�s�´������5�.4�Z~�U
����@�|&��~3�Ӽȉ�x׎e�5p��w���Э�P��~x�f`t8�u�|�@��gq����5$�|��vp�L ���5;�>�L	@ �)�u�
���]��������sJ�:7���L�U�`�a9�<y��O�� �A�3�{��TQ�v�u���ǌ�6yƏ��&vx�����	�cv>���(��&ĸ��"�I�2�[��Q�78{m���1W���K��U���'	��&L2IJ��-��2.M���5��W�?��J9�>\����o��8�m��yl��~�p�CCt�4�N���lT*,�c>X��a���T�� c{�K�-�x��_;�s�#�c*�P5r�q�����4#��z���%q�+,�1�mz�/�$?���"�w�B�ti<:BH� a���'�L�`�e�Pj�:�|ߧR(�`���~8�~:�N���a����'�ilH>�h)�3x�y�kM�������P,�Kd/
��� Rv1|����5���a¸V��97�L0��$	
�YOu�U��4B�c�և. 2&��r��U�nT=keBG*�h�M#�KU�⺄f�:��sL����{��&y.�ө��=ʒ��gO��q��X����PlB v*U�-1�*��.����BQ���r��?���r���>��"�!�}���(	�\w׻��j2"���.+뾹s�Z�Pu��(�֌�g���͘�0T�d>��%��iX8�x����n?�	�.%A��_|�1�k2ӹ1�	s(0#��v����횣��B�#JClx���!A�tt�<T�� -O�S8ɜ�t*Z@�?w	4
2$�v�����)�M`�-H�	��s��^W���"�>�^{/ʺ���`����p#��v�?O�Ť{�73�p
$5��JW�@ÔX� dӾ:H�\����w���A�4�#]pæ�	�M� ��R���p0�P.��u͐��u�������`{�4��2�y� �m�������IAXw>X �����z9X��;�Y�vZ�v���y<�����f���5�E�U*�X�p�N��h
b� �L����%3q�]I�bKgJ���Q��0������d��;��R,(֐���8<C��~�[�(�+�P���9�N��|�p��8H�B�,uL��\�I'b)e��� G&��X�7���C�}� ��Q���7��0���x4J�Ѓ�!�<
� "tCj�|g�ά�U�����I��"�p���&X�2!-3C��)(�qW9�������V��
>fwǍ:)�r��o�*�����|!�P��A{�񔂌7��~��@���_8k1�T��.�o��Ebi�Ty�FHn*L���/"XҠcY|��"^$��8����ĉi��^m�Ƌ� :n�mh��P�%
����,V���_i���:f�)D�� !;��c��k��"�>���b�&}n}<�"Lc;֦z�2���<����-�֏��6-����Ds(�$�fU���BXF�(g��Sr0@�q�7�I��-��n��,H;�<��$wȜx�ġ�R�L��Ԛ�
X`�����U�3�L ���̀:�m� �(a�|�ժ��ɓ���Q ��� ���L2W�J�΂���*�
����dX��URiWx&�P#$Vbh�O:���!�m{�rK�@�1�����w-X��7��>{㭀�'�voӳ��(�=\��b��~fp-E=�J)��˿�%# r-x�L-�VC�L�N
7�
Qm�c�1s�����Nb��sS�d�X����1�:��t:/U�*������&���>P��\S����F�`�{����L&��}oӆ"�:\qʸ=�XT����'�)�����»����Y�d9e��P9߱|c� y�D��1��<�	
ȧ�ǏW�ȩ�E��?o�tUZ�7/��+�4�X<fu�像4���le����sW�.�T��Ơ�SH��=f\�˗*�d��[��KQ�lΌc�:]�w<��?��q��{�p�8��Y�eϢOV�:{��P�.Qf�y����;�L!����������{�����x���]\�#��\� \�(�����H�L�>Y*)����|������?{2��&t�*8`0$��CSa�N�|�0,ȑn ���0�駧���b�`zv�.��HB~!��s?$�	NҦ�=vѱ�a�#��z<x}G�yg��QM�*/�K+�\~�D�s&v|R���i�y����G�kM}��<'�_�!zɊ^�u���|��{{���^��p��9��Lw�ՁP%[m@�m�V�D�6X*uq�o�Cа<�^�l���Vc�l��z��/-��j�wʡ�/����Ju�>2��FȀ޶�Xx���|F�?�T�?ף�1x���h�Zo����S#e����i��5��YGF���˖��#%Ms_�E2��^����z�,�����E�����ܒ�˲�EZ�PN�F���+!�@~����Ӟ��i��y�s�������%�/3�#�YV�6��%�����|����\�y��|�������Uض��R<e�5Z��)ay�%���ݸ\���j���d����~{��Ke���ƚ�����l�b֟��4�{T�!=�6kfr�8�(�:/��&�R�o�6�����Q��({�th��=��F�;(U��u��{bd�#�&'[~%��]
��N�pjn���ZA��iT��iA(!螱̷�/�JI�exMj��2xZװ��v|Y��ov�����IA�T4&1C^|���R7�?��-�9�A����D�lF���Ş7@�V��}-��L�2���⯵fb�*��m`N�gߎA��B(�����V����v����A�-����?N em�xبa%3_�OĂ�D��c=[���L��i�ɲ�&�	�n[����փ5oGPƏf�E�"ԅ��b%��Y��R��NCb�\sd�N15���MWx�&>o@q���f�ͿMCU�_ca��"(?��~�X��_��s��f���Y3o�D�����Xw��Ǣ�}9�Z�����L��*�|,�.�q��{c�5k@���s�Yk�H疜((!��w=�ì�0Z
bGJ�����*���4R=�RLޭ�R"Q2D�ԭ{_R�El]�1z��+:>׫K��|�n�����K}+��\Z{���p�n�;�j����G�u����^TGJS)*V�w?��1��LF����� [��/*T�1���NW2W�ˮ$���fǒ02em��%׫T"A�vОV���F�x��e��kl:�D�:���|�0����u�}d�y*��b�*��"�6���C��&�$}����H��h��O��|E��.<<�zD���b3���+�b*5u���	�hed���m��:Q�{p���+��YI�ֈ*d��V���h�kh>�\5�Bj��w7w���ʓ��'��+�s����FÖ�1c��-��l 	Z!���?����W�O7�>\�i�{O��^�7l+�y䔯U�� (#J�UO���x��=����k�:�J����qV�{.3��.[���"T�s&����X���e L��i�/~�Am;�M�{yр�����0���c�V�_�������9��]����`���� +��_�G��Ŵ�U�r�uA�_�G���.�BD���5�ފ�,�=�%���:XU�A�5��n ����ʀt��b�J�����D�n��o�mS�{z�������$1XCI	b��*/�d�G�px���1*rn���������\W��[� S��Jh��)���3Yx�#z�\R��v�G��Z08��^���yc:/O�O�o �K�#�{�(�&<*@ڟ����}t8��=+T��(�����ͧF�E�����>Z�@1�q�/k�o733G�HT�wqUX�ٻN����6��1��E�B���P���Y=�����e��g*=��BG�'�oE�X��s�����ZoB��@,�T_=�j)P���k�Xc���_LQ�'��Ih�|=�:��C���;l�%��_�IW�;�W�ǳd)��[��%:Pf�� JW����`]>H�J��3,i�L00��������g'@D����q��~�,;f�*P��Q���5%W@�/E�l0�ʢ�D(��1" }�:�u�A�����Ld��xhD)���_\��I!<Q��lc`*S|��{�e,;TX��Q��}�`ٳ�g��m��0J��drIB�@����vN'6͊�ݽ!r��F���f��Ο>��/u��c/$� �����Oׇ���cjm��"��ՊQ��~��o uG���]�j��%<Z��mK�T����h����OC�Ҧ�a�v~��
�.�3	�o]:�w+M���́'�
\�/�o ��>;>�R*���O:E���Φ&]�b�h�z1���y8�pxF�DŎ�f��B�$�^� ���>R���}���|جOֱ�Ӷ���p��=O���NY#6���^O��^� �t�̙���B�4�<��1`sœ;���*z�h��-�ɵ%A��a�VΔ�L���Y���xT-Z�¿M2>MH�YL|�q�+��>^��q�=ʌ�e���H2�)
#d�Fq0���&�	��4va�	�n�e%c�|#��i�w�@����X�{�w.��0� ;��Y�|���
��#�ᆅ�r!�r+�bv#P�69�i���� �Aڼ� ,� �P�1)Ui��匸TiH�8����2�\d�/dn �SNM �����d�jW�a𨟷��H&/q��t]ה�ϓ�%��B�@�B1dS
�T}�93�N�<�8��<M����������Sq^�Z����۟�z#eF|�S	x�3���8���O�N��q��
���t��uDW�3��-�����8�������b;���HЕ�r��9J���`,������Ap�����Sλ+ׅ�1[��Q�w�S>BJt�Jch��na�z9x�L��";���S\?�dm̽��w�Ǫ-��+L�yN��*��*Z��wjbdyE�;N$��Q-~��#���<���W�|�ɛ;;u!m����f#̗\���MU�$^�)=c�* �*�B��Cc��ކ�9�*T�lG���x5���G���z�e�=�����j2;*�%R�����{�H��%"���nFb�a�m��6�{!֮i�)�������?��7��q&�~��%���Ƿ���
�M%�fКv�
�l��4g�8�N�%�d�����H�W�A�%���0�$"�����l��'Tws����gݖ�yT���A��]�,dU�������,)���r~w����Б�W�
���g(��]��N2�`��/�q��
��*�Xķ���;��f�����"���ǲw�����|�&�(��k1�l��)H׃�%�$Y^f��%&�81qF��P�Z�vs\2��ɦ>v�!dn�w�{N�9�u�؋�_6��0�Q�N�ȷ$���5��s@�w�*��G�����=��-��<]|c���	���(����ScG� `�M{�rz\�;��l����_�;%�a�o$b���<�r��.�(����}�)���;O����lFҏx�[.��M$���r�C�M�΋�l�����)�CN	��aF�m�o䓾�ػ���xi�!PM#Ŏ��~޶�z1��m�j��Qo#[�Zp����\R4v�^���n;�m"^DI#�ĐD�֟�
��85s��m��ë�Ї����yVW:IR���Wc_7��Mc�㮙Nɕ���鹏F���y��P"1Rk[1\+�ϷwE� f2���Ī�yJ(��8�O`�_�	bf#:N���A��1����J5$��_�^g
���0�l�~�d��	}e�Q�k��;�W��#"�Es-�ܹv}�K3s�h��3�l�Բ�GN�Fn�^N��>e�Rp��ۦʈͨ��7Zz?��#�6�~�㹅C��W�i�N?�1|�9��Q �n��uh�f�${H��}#���v.<hk{n�Gg��&��o����?pw����'��O��I��9� ���j�M��C����a�.�"�p�i2���r}�r~�)9 �e���6��`������cP3d��6���Y�%VT8FВ��*�	��.�bV��h�hU�3�w��-���b�)��~�\c��VK%L/9<⚑�e��������df�����i	*C����N����~v6/�
�پ��;|�����9bE���+^���D2kĎb����V8��=��P����]���\Q򗁾��k�{�9~^c��(�M��mh�t�~6 �ob�1Z�R�A�o r��ic��(��gߖ�rE�l�{�(��:�dނcM�.%�y�����#�c� �����to��9�����.KS�-Y]�q�ҁx�=�˻��lY��޼ي����!�0�O��3��Ϋ�=�Z]�����'���b�2Ӓ��BԆ��lF�;� 
�f�A�ЋUʗՌ�2��m����9�#-ɰ�6���7N�1;`��
�K?���J��bT�����̂N]�(�����<\�5\ؿ�+b��c#�L�"�+��p	k��4q�?;�+�Q�\{

�+$3�鸛l�J	+ڴ3���w�cŏ9��y�����#z����Κ4��E�G�T����N�М#	��-R��ĥ g�ԃ��l�n٘d$�B	~z6��@�@�.#����o�V|���%c��Q�����V�^��|�oGK���+�G8;�����^�A���v�$�Ԏg�i�������6ꊾ�XlYo�ӡs�b�m_�#�_�q��}}b�Q�0���}[��1�	翄e)%�z4/�anɠ��j�K07:�yZ՚0�� �bɇ�F�y�!�I配$��c��ps���@����U_�b����#�9$Я�#��L`�υ�����lbA`�l�:��#�%����\.������ja硩g3�:����L"Wt�al�H�>un�Ș�_�tY���G�{� A#Ow��D-mH>�i Oʜpc#}I3eqLn6��QMD2����]�5͊E����(�7�nk�7C�
u��e�?3���A��Z��/2u,	�t��U	Vtty�_�g′�V3U�Z�-�i��ȿ���!Ngq��!��S� 'ҩ��Ȍt5�z�$�U8�.M�����Ā�)��TL�Om�On疒:�����j�h��s!�ۨ� d�_A{�#y�ʆ6l��{9BT��bIi�ٰ��� +Zg��=:�����¿�-��dm���=�Z� �P$�[��OH�T7���(������q�<�$t�����]nu��%%5�=s�R����G(R��f���b9�ỻ�<�M1�����{+^?�m�)�r�)�T�|��9�����U����V޹���)��1����Y|�Ǜ<�2~�@�z��L��2�w��y5�).ma~F��a�D5�g����Ě�e�Ԛ��@M� �*gc/E�tq�YT��c�Xl���wU��a��B%x��萐����A Gݡz����Y�_>~�@e7�����=�[s�}}�(p��/h��8)�\��mޟ$m�U�k_%�,HjAغN��):��B�P�=�;� 8~!�LEھ��ߍϩx�D�򦿁Cg�M�Q�gZ&po�p�/��l�U0��E !+6p��(�:)�@/�,)�yUzi+H���O��	_o[�@T:��1��ǶQ�V�3J0v��u��)@
�o!/����ȚI�fE��~6��<�>c6�Ou�n�{��������ŏ��
�lz�SQ()��ۜ93P�Q����i�2��T��5qE���F��U�"����
�"<�`�iC]_�EKi��2����R/��9��O�cDѝ�3e���p��7��_��hjNL��Xh�a���M�1�D�2�D�O��we�CqO�[��އ�����9�����)qnlX��N�I]"�1��Ҟ/�:bR�댆 C=�P�Aw��;��XFK������#6��sG[���G2'R-%�|r���\�����CIm�����U2#��g%m+_�8�~��be�����!d��eo�,:*ߙW�%B�\��&��{�䳧���	!!�����?^��G����E�f}Y{	V��)�E�����D�-��]4�u8-�EKP8��&q�^�.�h�?w�x�ۏ y�Љ�}�iy��H3�c����zɱZ�@Jm�j1v�Vb"��ϵI�1��3������ �X�G�G�V�{O&�^Җ"|��U8&h��U5&��[�B:d�Y�3�k�Eu�R|	"��*�����J�v�����!��X�%������	�C�U�tF���C�^�BB1h�  7�ݴ60+Y������b�d�fbr�TҐQK��y��q�2����6E[d���z�0�V6)��'tS����9Xo �r����e�=,�)������_��[sO+y��f+���sw�ye=Q,�=�����Ů���@ź���J��c�S���4 ���|�ߔ���`��o���J��I���w��4���|vt�4����s�$WB�$ߕ*ȃ����@��lp@�B�p�%���b�ϟ�N��N��s;��Y��J���ڛ'�⦭�K���樻���Kʆ5�ܐՌ�}��i����/�O��#�wʮ�O���C��٣��ޅ���g`mi�u���eʳY��rq>ϋ�~@���q睻���n0T�ՔJ]C|������zϟ-�r,�_+.:?�ͣ�m>༚Dh��)�ݵ/�WG��w��<���I���"�����}_ZV�y/�3���5o[,����<mm���������ja���:���1Nɠ|0Ws�:Wk���ѽ���s��c��@�O�[�(s9f+�֒��U�Ȼ����@��R_)E���sE�UgAGǓ�J���;�dW�4�B>����!-��[f���u�j��H���{���2�9m�em�׋�A5S�Ć�F���kq���T��'����p[�`�M9f�H��w%��	B�A�Q�=)�O��0������5����Ww��v1t����W;=;�	�Su=4%��y}4���r�>Ų����N@'G��5��x�#�r+ ��4�
��\��9�"��*�~�&_;JB:�rR���xH;q�Ó<�c؅�fP�a��_��MccpQXT	_@M~��j�
� �9�@�~��\�*�ۤ�iLnk�.�pLyux/��e�;�4�~�����l���;��'$y�&J��"�c,��^
t�Bcs�-��$�����8H~q�+W���_H+����m�h��.]S�Q@�v+�Ʃ��|�jA���c����*���.V� 3=�ڈ�p�ݔ8��]|n��(��i�-B)���>�<cg޸�X�:�����������襝�\�L���~DW#�=Y��:.���J2���!>�D%�O�U.c��YB�%o�:4��qpa����$����Li� ��r`���j3�5W�l��tGS���_+��>KR�!��$_U��0��^�Y��w����!���e���8�Qi����>)N�[�;L�v�D� 
m�JLFx̢��H��q�5>���1z��᫥�|�	)��K�5ԑ'E7�5�p�T��Y y��;������[�N��e�Iq�%�6VR�@l�*  .�=���7 MaI�`�n���}>�f7����hz�:,a?�l�����hw0��M�Y�HU���U=#J�it9�3�ڠ���.�ҏ��X{Z�������E�Eg��rb�5�4��Sno�����PU+X�LmqMk���՗�풍�	��Ġ��X�-��絞K	O�{�Q7�/�i����6��,��K
r����[�>9����/����]��A=hTi ��r��qw+�v��w��KD�'���g1����h8#0��F�	��k�
k�D��x��ܧ�+�3L�]-�t}��`����]W|��VV��Ҳ�抟?���+}ٴ@u������ �';�1�li���	�]��������t,��Yj>v妉Ng�Y��H.	�}N�UW���xu��D y���V�b�F�aC�G��A"Oăܛp!������0[����ӻ,y$b�˄���`?�#6ܦ��$��o!�3 �D��襭@�_�Ы��Q��|~lw�/�i �?��y!35�=�:���PL>S�='d�$P�� ������s��y�i��tT��ae���*���u��R�#�R�����q�VDo]�ڃz+n f��
��	�A�0O�/��.��q���ъ �-�_=�'��ڽZ�e� %�7��w��y��yb�1��~h�u���&J���iA7@j��V�<������,�PK   �rUh�NS  #     jsons/user_defined.json��]K�0����u�~��-�@�8�F��#��.�I���ݓ�9a]�r��>�'9;�m[�b�k�^*Vs�*d��4�L����H5��w��"_�mê	�Q0�N	�2��J�-H�#p'�7���0�˚8Է=B��Q������:�7u����t�Ɲ��w���R�#����x�֮��r1�D��~�r�6�6���"uAul�ˍiQ�`��0�I/�{	ļZv���y<#����7���빘�	�(���L��L��R��0i������xz�����y���Y�s��/�/��|��\�Ogh����0��+X�JJ�Lu|��f�J).ܐ!>PK   �rUB/  �c             ��    cirkitFile.jsonPK   �rU�#��g (t /           ��\  images/85cf0215-4010-4105-9e1b-ea712a483bd2.jpgPK   �rUh�NS  #             ��3s jsons/user_defined.jsonPK      �   �t   